

    module v$ROM1_462(q, a, clk);
    output reg [0:0] q;
    input clk;
    input [11:0] a;
    reg [0:0] rom [4095:0];
    always @(posedge clk) q <= rom[a];
    integer i;
    initial
    begin
        for (i=0; i < 4096; i=i+1)
        begin
            rom[i] = 0;
        end
        q = 0;
    
        rom[0] = 0;
rom[1] = 1;
rom[2] = 0;
rom[3] = 0;
rom[4] = 0;
rom[5] = 1;
rom[6] = 0;
rom[7] = 0;
rom[8] = 0;
rom[9] = 1;
rom[10] = 1;
rom[11] = 1;
rom[12] = 0;
rom[13] = 0;
rom[14] = 1;
rom[15] = 0;
rom[16] = 0;
rom[17] = 0;
rom[18] = 0;
rom[19] = 0;
rom[20] = 0;
rom[21] = 1;
rom[22] = 1;
rom[23] = 1;
rom[24] = 1;
rom[25] = 0;
rom[26] = 0;
rom[27] = 0;
rom[28] = 0;
rom[29] = 0;
rom[30] = 0;
rom[31] = 1;
rom[32] = 1;
rom[33] = 1;
rom[34] = 1;
rom[35] = 1;
rom[36] = 1;
rom[37] = 1;
rom[38] = 1;
rom[39] = 1;
rom[40] = 1;
rom[41] = 1;
rom[42] = 1;
rom[43] = 1;
rom[44] = 1;
rom[45] = 1;
rom[46] = 1;
rom[47] = 1;
rom[48] = 1;
rom[49] = 1;
rom[50] = 1;
rom[51] = 1;
rom[52] = 1;
rom[53] = 1;
rom[54] = 1;
rom[55] = 1;
rom[56] = 1;
rom[57] = 1;
rom[58] = 1;
rom[59] = 1;
rom[60] = 1;
rom[61] = 1;
rom[62] = 1;
rom[63] = 1;
rom[64] = 1;
rom[65] = 1;
rom[66] = 1;
rom[67] = 1;
rom[68] = 1;
rom[69] = 1;
rom[70] = 1;
rom[71] = 1;
rom[72] = 1;
rom[73] = 1;
rom[74] = 1;
rom[75] = 1;
rom[76] = 1;
rom[77] = 1;
rom[78] = 1;
rom[79] = 1;
rom[80] = 1;
rom[81] = 1;
rom[82] = 1;
rom[83] = 1;
rom[84] = 1;
rom[85] = 1;
rom[86] = 1;
rom[87] = 1;
rom[88] = 1;
rom[89] = 1;
rom[90] = 1;
rom[91] = 1;
rom[92] = 1;
rom[93] = 1;
rom[94] = 1;
rom[95] = 1;
    end
    endmodule
     

    module v$RAM0_1680(q, a, d, we, clk);
    output reg [15:0] q;
    input [15:0] d;
    input [11:0] a;
    input we, clk;
    reg [15:0] ram [4095:0];
     always @(posedge clk) begin
         if (we)
             ram[a] <= d;
         q <= ram[a];
     end

    integer i;
    initial
    begin
        for (i=0; i < 4096; i=i+1)
        begin
            ram[i] = 0;
        end

        q = 0;

        ram[0] = 8192;
ram[1] = 838;
ram[2] = 1862;
ram[3] = 32769;
ram[4] = 1862;
ram[5] = 32769;
ram[6] = 322;
ram[7] = 28672;
ram[2036] = 50786;
ram[2037] = 205;
ram[2038] = 3281;
ram[2039] = 12997;
ram[2040] = 3797;
ram[2041] = 35840;
ram[2042] = 15561;
ram[2043] = 3285;
ram[2044] = 717;
ram[2045] = 3793;
ram[2046] = 50688;
    end
    endmodule

    

    module v$data$ram_1818(q, a, d, we, clk);
    output reg [15:0] q;
    input [15:0] d;
    input [11:0] a;
    input we, clk;
    reg [15:0] ram [4095:0];
     always @(posedge clk) begin
         if (we)
             ram[a] <= d;
         q <= ram[a];
     end

    integer i;
    initial
    begin
        for (i=0; i < 4096; i=i+1)
        begin
            ram[i] = 0;
        end

        q = 0;

        ram[0] = 15360;
ram[1] = 14336;
ram[2] = 12629;
ram[3] = 65535;
ram[4] = 8260;
ram[5] = 13312;
ram[6] = 85;
ram[7] = 0;
    end
    endmodule

    

    module v$RAM1_13398(q, a, d, we, clk);
    output reg [15:0] q;
    input [15:0] d;
    input [11:0] a;
    input we, clk;
    reg [15:0] ram [4095:0];
     always @(posedge clk) begin
         if (we)
             ram[a] <= d;
         q <= ram[a];
     end

    integer i;
    initial
    begin
        for (i=0; i < 4096; i=i+1)
        begin
            ram[i] = 0;
        end

        q = 0;

        ram[0] = 8192;
ram[1] = 722;
ram[2] = 3798;
ram[3] = 0;
ram[4] = 0;
ram[5] = 0;
ram[6] = 0;
ram[7] = 1742;
ram[8] = 32769;
ram[9] = 4099;
ram[10] = 28672;
ram[2036] = 50786;
ram[2037] = 205;
ram[2038] = 3281;
ram[2039] = 12997;
ram[2040] = 3797;
ram[2041] = 35840;
ram[2042] = 15561;
ram[2043] = 3285;
ram[2044] = 717;
ram[2045] = 3793;
ram[2046] = 50688;
    end
    endmodule

    
module main (
	clk,
	v$DIV$INST0_6905_out0,
	v$DIV$INST1_7011_out0,
	v$IR1_6873_out0,
	v$BYTE$RECEIVED_11192_out0,
	v$IR0_13305_out0,
	v$R13_375_out0,
	v$R11_398_out0,
	v$R00_3807_out0,
	v$R02_6966_out0,
	v$R12_10714_out0,
	v$R10_11216_out0,
	v$R03_13304_out0,
	v$R01_13752_out0,
	v$REGISTER$INUP16_384_out0,
	v$REGISTER$INUP0_12240_out0,
	v$REGISTER14_3201_out0,
	v$REGISTER15_8833_out0);
input clk;
input v$DIV$INST0_6905_out0;
input v$DIV$INST1_7011_out0;
output  [11:0] v$REGISTER14_3201_out0;
output  [11:0] v$REGISTER15_8833_out0;
output  [15:0] v$IR0_13305_out0;
output  [15:0] v$IR1_6873_out0;
output  [15:0] v$R00_3807_out0;
output  [15:0] v$R01_13752_out0;
output  [15:0] v$R02_6966_out0;
output  [15:0] v$R03_13304_out0;
output  [15:0] v$R10_11216_out0;
output  [15:0] v$R11_398_out0;
output  [15:0] v$R12_10714_out0;
output  [15:0] v$R13_375_out0;
output  [15:0] v$REGISTER$INUP0_12240_out0;
output  [15:0] v$REGISTER$INUP16_384_out0;
output  [7:0] v$BYTE$RECEIVED_11192_out0;
reg  [11:0] v$REG1_432_out0 = 12'h0;
reg  [11:0] v$REG1_433_out0 = 12'h0;
reg  [11:0] v$REG1_7134_out0 = 12'h0;
reg  [15:0] v$IHOLD$REGISTER_2013_out0 = 16'h0;
reg  [15:0] v$IHOLD$REGISTER_2014_out0 = 16'h0;
reg  [15:0] v$REG0_10912_out0 = 16'h0;
reg  [15:0] v$REG0_10913_out0 = 16'h0;
reg  [15:0] v$REG1_13338_out0 = 16'h0;
reg  [15:0] v$REG1_13339_out0 = 16'h0;
reg  [15:0] v$REG1_2314_out0 = 16'h0;
reg  [15:0] v$REG1_2315_out0 = 16'h0;
reg  [15:0] v$REG2_12251_out0 = 16'h0;
reg  [15:0] v$REG2_12252_out0 = 16'h0;
reg  [15:0] v$REG3_4747_out0 = 16'h0;
reg  [15:0] v$REG3_4748_out0 = 16'h0;
reg  [1:0] v$REG1_10368_out0 = 2'h0;
reg  [1:0] v$REG1_7031_out0 = 2'h0;
reg  [7:0] v$REG1_10546_out0 = 8'h0;
reg  [7:0] v$REG1_2677_out0 = 8'h0;
reg v$FF1_10325_out0 = 1'b0;
reg v$FF1_10326_out0 = 1'b0;
reg v$FF1_13511_out0 = 1'b0;
reg v$FF1_1955_out0 = 1'b0;
reg v$FF1_4717_out0 = 1'b0;
reg v$FF1_4718_out0 = 1'b0;
reg v$FF1_4719_out0 = 1'b0;
reg v$FF1_4720_out0 = 1'b0;
reg v$FF1_4721_out0 = 1'b0;
reg v$FF1_4722_out0 = 1'b0;
reg v$FF1_4723_out0 = 1'b0;
reg v$FF1_4724_out0 = 1'b0;
reg v$FF1_4725_out0 = 1'b0;
reg v$FF1_4726_out0 = 1'b0;
reg v$FF1_4727_out0 = 1'b0;
reg v$FF1_4728_out0 = 1'b0;
reg v$FF1_4729_out0 = 1'b0;
reg v$FF1_4730_out0 = 1'b0;
reg v$FF1_4731_out0 = 1'b0;
reg v$FF1_4732_out0 = 1'b0;
reg v$FF1_4841_out0 = 1'b0;
reg v$FF1_48_out0 = 1'b0;
reg v$FF1_49_out0 = 1'b0;
reg v$FF2_11062_out0 = 1'b0;
reg v$FF2_2833_out0 = 1'b0;
reg v$FF3_11046_out0 = 1'b0;
reg v$FF3_2016_out0 = 1'b0;
reg v$FF3_2017_out0 = 1'b0;
reg v$FF4_2106_out0 = 1'b0;
reg v$FF4_2107_out0 = 1'b0;
reg v$FF4_463_out0 = 1'b0;
reg v$FF5_7100_out0 = 1'b0;
reg v$FF6_112_out0 = 1'b0;
reg v$FF7_2670_out0 = 1'b0;
reg v$FF7_2671_out0 = 1'b0;
reg v$FF7_2672_out0 = 1'b0;
reg v$FF7_2673_out0 = 1'b0;
reg v$FF7_4781_out0 = 1'b0;
reg v$FF8_10849_out0 = 1'b0;
reg v$FF8_10850_out0 = 1'b0;
reg v$FF8_10851_out0 = 1'b0;
reg v$FF8_10852_out0 = 1'b0;
reg v$FF8_11222_out0 = 1'b0;
reg v$FF9_8805_out0 = 1'b0;
reg v$REG1_11130_out0 = 1'b0;
reg v$REG1_11131_out0 = 1'b0;
wire  [10:0] v$C1_606_out0;
wire  [10:0] v$C1_607_out0;
wire  [10:0] v$C_1807_out0;
wire  [10:0] v$C_1808_out0;
wire  [10:0] v$IN1_10992_out0;
wire  [10:0] v$IN1_10993_out0;
wire  [10:0] v$IN1_13711_out0;
wire  [10:0] v$IN1_13712_out0;
wire  [10:0] v$IN1_2189_out0;
wire  [10:0] v$IN1_2190_out0;
wire  [10:0] v$IN1_2848_out0;
wire  [10:0] v$IN1_2849_out0;
wire  [10:0] v$IN_13668_out0;
wire  [10:0] v$IN_13669_out0;
wire  [10:0] v$MUX1_2401_out0;
wire  [10:0] v$MUX1_2402_out0;
wire  [10:0] v$MUX1_7143_out0;
wire  [10:0] v$MUX1_7144_out0;
wire  [10:0] v$MUX1_7702_out0;
wire  [10:0] v$MUX1_7703_out0;
wire  [10:0] v$MUX2_188_out0;
wire  [10:0] v$MUX2_189_out0;
wire  [10:0] v$MUX3_13312_out0;
wire  [10:0] v$MUX3_13313_out0;
wire  [10:0] v$MUX4_552_out0;
wire  [10:0] v$MUX4_553_out0;
wire  [10:0] v$MUX5_13670_out0;
wire  [10:0] v$MUX5_13671_out0;
wire  [10:0] v$OP2$SIG$NEW_11190_out0;
wire  [10:0] v$OP2$SIG$NEW_11191_out0;
wire  [10:0] v$OP2$SIG$NEW_11218_out0;
wire  [10:0] v$OP2$SIG$NEW_11219_out0;
wire  [10:0] v$OP2$SIG11_14_out0;
wire  [10:0] v$OP2$SIG11_15_out0;
wire  [10:0] v$OP2$SIG11_4827_out0;
wire  [10:0] v$OP2$SIG11_4828_out0;
wire  [10:0] v$OP2$SIG_13314_out0;
wire  [10:0] v$OP2$SIG_13315_out0;
wire  [10:0] v$OUT1_1873_out0;
wire  [10:0] v$OUT1_1874_out0;
wire  [10:0] v$OUT1_1972_out0;
wire  [10:0] v$OUT1_1973_out0;
wire  [10:0] v$OUT1_3294_out0;
wire  [10:0] v$OUT1_3295_out0;
wire  [10:0] v$OUT1_3853_out0;
wire  [10:0] v$OUT1_3854_out0;
wire  [10:0] v$Q_10339_out0;
wire  [10:0] v$Q_10340_out0;
wire  [10:0] v$Q_10341_out0;
wire  [10:0] v$Q_10342_out0;
wire  [10:0] v$RD$SIG$NEW_10872_out0;
wire  [10:0] v$RD$SIG$NEW_10873_out0;
wire  [10:0] v$RD$SIG$NEW_8759_out0;
wire  [10:0] v$RD$SIG$NEW_8760_out0;
wire  [10:0] v$RD$SIG11_7132_out0;
wire  [10:0] v$RD$SIG11_7133_out0;
wire  [10:0] v$RD$SIG11_8854_out0;
wire  [10:0] v$RD$SIG11_8855_out0;
wire  [10:0] v$RD$SIG_109_out0;
wire  [10:0] v$RD$SIG_110_out0;
wire  [10:0] v$SEL2_13496_out0;
wire  [10:0] v$SEL2_13497_out0;
wire  [10:0] v$SHIFTED$SIG_10802_out0;
wire  [10:0] v$SHIFTED$SIG_10803_out0;
wire  [10:0] v$SHIFTED$SIG_13632_out0;
wire  [10:0] v$SHIFTED$SIG_13633_out0;
wire  [10:0] v$SIG$RD$11bit_3301_out0;
wire  [10:0] v$SIG$RD$11bit_3302_out0;
wire  [10:0] v$SIG$RM$11bit_6892_out0;
wire  [10:0] v$SIG$RM$11bit_6893_out0;
wire  [10:0] v$SIG$TO$SHIFT_10712_out0;
wire  [10:0] v$SIG$TO$SHIFT_10713_out0;
wire  [10:0] v$SIG$TO$SHIFT_5836_out0;
wire  [10:0] v$SIG$TO$SHIFT_5837_out0;
wire  [10:0] v$_13310_out0;
wire  [10:0] v$_13311_out0;
wire  [10:0] v$_13484_out0;
wire  [10:0] v$_13485_out0;
wire  [10:0] v$_13761_out0;
wire  [10:0] v$_13762_out0;
wire  [10:0] v$_2026_out0;
wire  [10:0] v$_2027_out0;
wire  [10:0] v$_2028_out0;
wire  [10:0] v$_2029_out0;
wire  [10:0] v$_2030_out0;
wire  [10:0] v$_2031_out0;
wire  [10:0] v$_2032_out0;
wire  [10:0] v$_2033_out0;
wire  [10:0] v$_2034_out0;
wire  [10:0] v$_2035_out0;
wire  [10:0] v$_2036_out0;
wire  [10:0] v$_2037_out0;
wire  [10:0] v$_2038_out0;
wire  [10:0] v$_2039_out0;
wire  [10:0] v$_2040_out0;
wire  [10:0] v$_2041_out0;
wire  [10:0] v$_2042_out0;
wire  [10:0] v$_2043_out0;
wire  [10:0] v$_2044_out0;
wire  [10:0] v$_2045_out0;
wire  [10:0] v$_2046_out0;
wire  [10:0] v$_2047_out0;
wire  [10:0] v$_2048_out0;
wire  [10:0] v$_2049_out0;
wire  [10:0] v$_2050_out0;
wire  [10:0] v$_2051_out0;
wire  [10:0] v$_2052_out0;
wire  [10:0] v$_2053_out0;
wire  [10:0] v$_2054_out0;
wire  [10:0] v$_2055_out0;
wire  [10:0] v$_2191_out0;
wire  [10:0] v$_2192_out0;
wire  [10:0] v$_2771_out0;
wire  [10:0] v$_2772_out0;
wire  [10:0] v$_2834_out0;
wire  [10:0] v$_2835_out0;
wire  [10:0] v$_2836_out0;
wire  [10:0] v$_2837_out0;
wire  [10:0] v$_2971_out0;
wire  [10:0] v$_2972_out0;
wire  [10:0] v$_4591_out0;
wire  [10:0] v$_4592_out0;
wire  [10:0] v$_4733_out0;
wire  [10:0] v$_4734_out0;
wire  [10:0] v$_7714_out0;
wire  [10:0] v$_7715_out0;
wire  [10:0] v$shifted1_2666_out0;
wire  [10:0] v$shifted1_2667_out0;
wire  [11:0] v$A1_11043_out0;
wire  [11:0] v$A1_7019_out0;
wire  [11:0] v$A1_7020_out0;
wire  [11:0] v$ADDER$IN_10995_out0;
wire  [11:0] v$ADDER$IN_10996_out0;
wire  [11:0] v$ADDRESS0_10982_out0;
wire  [11:0] v$ADDRESS1_2854_out0;
wire  [11:0] v$ADDRESS_4662_out0;
wire  [11:0] v$ADRESS$ins0_11169_out0;
wire  [11:0] v$ADRESS$ins1_10617_out0;
wire  [11:0] v$ADRESS0_11217_out0;
wire  [11:0] v$ADRESS1_1906_out0;
wire  [11:0] v$ADRESS_2339_out0;
wire  [11:0] v$ADRESS_2340_out0;
wire  [11:0] v$ADRESS_2542_out0;
wire  [11:0] v$ADRESS_2543_out0;
wire  [11:0] v$ADRESS_8683_out0;
wire  [11:0] v$A_10821_out0;
wire  [11:0] v$A_10822_out0;
wire  [11:0] v$C1_2426_out0;
wire  [11:0] v$C1_2427_out0;
wire  [11:0] v$C1_3210_out0;
wire  [11:0] v$C1_3211_out0;
wire  [11:0] v$C2_10761_out0;
wire  [11:0] v$C2_10762_out0;
wire  [11:0] v$C2_2413_out0;
wire  [11:0] v$EA_13516_out0;
wire  [11:0] v$EA_13517_out0;
wire  [11:0] v$JUMPADRESS_4745_out0;
wire  [11:0] v$JUMPADRESS_4746_out0;
wire  [11:0] v$JUMPADRESS_6964_out0;
wire  [11:0] v$JUMPADRESS_6965_out0;
wire  [11:0] v$MULTI$PRODUCT_7104_out0;
wire  [11:0] v$MULTI$PRODUCT_7105_out0;
wire  [11:0] v$MUX1_10773_out0;
wire  [11:0] v$MUX1_10774_out0;
wire  [11:0] v$MUX1_7097_out0;
wire  [11:0] v$MUX2_13656_out0;
wire  [11:0] v$MUX2_13657_out0;
wire  [11:0] v$MUX3_10330_out0;
wire  [11:0] v$MUX3_10331_out0;
wire  [11:0] v$MUX3_3225_out0;
wire  [11:0] v$MUX3_3226_out0;
wire  [11:0] v$MUX4_2658_out0;
wire  [11:0] v$MUX4_2659_out0;
wire  [11:0] v$MUX5_10845_out0;
wire  [11:0] v$MUX5_10846_out0;
wire  [11:0] v$MUX8_13785_out0;
wire  [11:0] v$MUX8_13786_out0;
wire  [11:0] v$NEXT$ADRESS_3243_out0;
wire  [11:0] v$NEXT$ADRESS_3244_out0;
wire  [11:0] v$NEXTADD_10526_out0;
wire  [11:0] v$NEXTADD_10527_out0;
wire  [11:0] v$NEXTADRESS_1803_out0;
wire  [11:0] v$NEXTADRESS_1804_out0;
wire  [11:0] v$NOUSED_13492_out0;
wire  [11:0] v$NOUSED_13493_out0;
wire  [11:0] v$PC$COUNTER$NEXT_7064_out0;
wire  [11:0] v$PC$COUNTER$NEXT_7065_out0;
wire  [11:0] v$PC$COUNTER_25_out0;
wire  [11:0] v$PC$COUNTER_26_out0;
wire  [11:0] v$RAM$ADDRES$MUX_13649_out0;
wire  [11:0] v$RAM$ADDRES$MUX_13650_out0;
wire  [11:0] v$RAM$ADDRESS$MUX_8803_out0;
wire  [11:0] v$RAM$ADDRESS$MUX_8804_out0;
wire  [11:0] v$RAMADDRMUX_10542_out0;
wire  [11:0] v$RAMADDRMUX_10543_out0;
wire  [11:0] v$RAMADDRMUX_2232_out0;
wire  [11:0] v$RAMADDRMUX_2233_out0;
wire  [11:0] v$RAMADDRMUX_7066_out0;
wire  [11:0] v$RAMADDRMUX_7067_out0;
wire  [11:0] v$RAMADDRMUX_92_out0;
wire  [11:0] v$RAMADDRMUX_93_out0;
wire  [11:0] v$REGISTER4_1705_out0;
wire  [11:0] v$REGISTER4_1706_out0;
wire  [11:0] v$REGISTER_13346_out0;
wire  [11:0] v$REGISTER_13347_out0;
wire  [11:0] v$REGISTER_216_out0;
wire  [11:0] v$REGISTER_217_out0;
wire  [11:0] v$SEL7_4850_out0;
wire  [11:0] v$SEL7_4851_out0;
wire  [11:0] v$SEL8_10686_out0;
wire  [11:0] v$SEL8_10687_out0;
wire  [11:0] v$_10370_out0;
wire  [11:0] v$_10371_out0;
wire  [11:0] v$_10783_out0;
wire  [11:0] v$_10784_out0;
wire  [11:0] v$_107_out0;
wire  [11:0] v$_108_out0;
wire  [11:0] v$_11137_out0;
wire  [11:0] v$_11138_out0;
wire  [11:0] v$_11139_out0;
wire  [11:0] v$_11140_out0;
wire  [11:0] v$_13291_out1;
wire  [11:0] v$_13292_out1;
wire  [11:0] v$_224_out0;
wire  [11:0] v$_225_out0;
wire  [11:0] v$_2411_out0;
wire  [11:0] v$_2412_out0;
wire  [11:0] v$_2439_out0;
wire  [11:0] v$_2440_out0;
wire  [11:0] v$_2793_out0;
wire  [11:0] v$_2794_out0;
wire  [11:0] v$_2795_out0;
wire  [11:0] v$_2796_out0;
wire  [11:0] v$_2797_out0;
wire  [11:0] v$_2798_out0;
wire  [11:0] v$_2799_out0;
wire  [11:0] v$_2800_out0;
wire  [11:0] v$_2801_out0;
wire  [11:0] v$_2802_out0;
wire  [11:0] v$_2803_out0;
wire  [11:0] v$_2804_out0;
wire  [11:0] v$_2805_out0;
wire  [11:0] v$_2806_out0;
wire  [11:0] v$_2807_out0;
wire  [11:0] v$_2808_out0;
wire  [11:0] v$_2809_out0;
wire  [11:0] v$_2810_out0;
wire  [11:0] v$_2811_out0;
wire  [11:0] v$_2812_out0;
wire  [11:0] v$_2813_out0;
wire  [11:0] v$_2814_out0;
wire  [11:0] v$_2815_out0;
wire  [11:0] v$_2816_out0;
wire  [11:0] v$_2817_out0;
wire  [11:0] v$_2818_out0;
wire  [11:0] v$_2819_out0;
wire  [11:0] v$_2820_out0;
wire  [11:0] v$_2821_out0;
wire  [11:0] v$_2822_out0;
wire  [11:0] v$_3035_out0;
wire  [11:0] v$_3036_out0;
wire  [11:0] v$_4488_out1;
wire  [11:0] v$_4489_out1;
wire  [11:0] v$_4585_out1;
wire  [11:0] v$_4586_out1;
wire  [11:0] v$_5846_out0;
wire  [11:0] v$_5847_out0;
wire  [11:0] v$_7116_out0;
wire  [11:0] v$_7117_out0;
wire  [12:0] v$_164_out0;
wire  [12:0] v$_165_out0;
wire  [12:0] v$_1825_out0;
wire  [12:0] v$_1826_out0;
wire  [12:0] v$_1827_out0;
wire  [12:0] v$_1828_out0;
wire  [12:0] v$_1829_out0;
wire  [12:0] v$_1830_out0;
wire  [12:0] v$_1831_out0;
wire  [12:0] v$_1832_out0;
wire  [12:0] v$_1833_out0;
wire  [12:0] v$_1834_out0;
wire  [12:0] v$_1835_out0;
wire  [12:0] v$_1836_out0;
wire  [12:0] v$_1837_out0;
wire  [12:0] v$_1838_out0;
wire  [12:0] v$_1839_out0;
wire  [12:0] v$_1840_out0;
wire  [12:0] v$_1841_out0;
wire  [12:0] v$_1842_out0;
wire  [12:0] v$_1843_out0;
wire  [12:0] v$_1844_out0;
wire  [12:0] v$_1845_out0;
wire  [12:0] v$_1846_out0;
wire  [12:0] v$_1847_out0;
wire  [12:0] v$_1848_out0;
wire  [12:0] v$_1849_out0;
wire  [12:0] v$_1850_out0;
wire  [12:0] v$_1851_out0;
wire  [12:0] v$_1852_out0;
wire  [12:0] v$_1853_out0;
wire  [12:0] v$_1854_out0;
wire  [12:0] v$_3192_out0;
wire  [12:0] v$_3193_out0;
wire  [12:0] v$_3194_out0;
wire  [12:0] v$_3195_out0;
wire  [12:0] v$_5851_out0;
wire  [12:0] v$_5852_out0;
wire  [12:0] v$_9802_out0;
wire  [12:0] v$_9803_out0;
wire  [13:0] v$_10767_out0;
wire  [13:0] v$_10768_out0;
wire  [13:0] v$_11049_out0;
wire  [13:0] v$_11050_out0;
wire  [13:0] v$_11055_out0;
wire  [13:0] v$_11056_out0;
wire  [13:0] v$_173_out0;
wire  [13:0] v$_174_out0;
wire  [13:0] v$_175_out0;
wire  [13:0] v$_176_out0;
wire  [13:0] v$_4483_out1;
wire  [13:0] v$_4484_out1;
wire  [13:0] v$_4549_out0;
wire  [13:0] v$_4550_out0;
wire  [13:0] v$_4551_out0;
wire  [13:0] v$_4552_out0;
wire  [13:0] v$_4553_out0;
wire  [13:0] v$_4554_out0;
wire  [13:0] v$_4555_out0;
wire  [13:0] v$_4556_out0;
wire  [13:0] v$_4557_out0;
wire  [13:0] v$_4558_out0;
wire  [13:0] v$_4559_out0;
wire  [13:0] v$_4560_out0;
wire  [13:0] v$_4561_out0;
wire  [13:0] v$_4562_out0;
wire  [13:0] v$_4563_out0;
wire  [13:0] v$_4564_out0;
wire  [13:0] v$_4565_out0;
wire  [13:0] v$_4566_out0;
wire  [13:0] v$_4567_out0;
wire  [13:0] v$_4568_out0;
wire  [13:0] v$_4569_out0;
wire  [13:0] v$_4570_out0;
wire  [13:0] v$_4571_out0;
wire  [13:0] v$_4572_out0;
wire  [13:0] v$_4573_out0;
wire  [13:0] v$_4574_out0;
wire  [13:0] v$_4575_out0;
wire  [13:0] v$_4576_out0;
wire  [13:0] v$_4577_out0;
wire  [13:0] v$_4578_out0;
wire  [13:0] v$_4816_out1;
wire  [13:0] v$_4817_out1;
wire  [13:0] v$_538_out0;
wire  [13:0] v$_539_out0;
wire  [13:0] v$_627_out1;
wire  [13:0] v$_628_out1;
wire  [14:0] v$CIN_2356_out0;
wire  [14:0] v$CIN_2371_out0;
wire  [14:0] v$REST_162_out0;
wire  [14:0] v$REST_163_out0;
wire  [14:0] v$_10354_out0;
wire  [14:0] v$_10355_out0;
wire  [14:0] v$_10455_out0;
wire  [14:0] v$_10456_out0;
wire  [14:0] v$_10457_out0;
wire  [14:0] v$_10458_out0;
wire  [14:0] v$_10651_out0;
wire  [14:0] v$_10652_out0;
wire  [14:0] v$_10653_out0;
wire  [14:0] v$_10654_out0;
wire  [14:0] v$_10655_out0;
wire  [14:0] v$_10656_out0;
wire  [14:0] v$_10657_out0;
wire  [14:0] v$_10658_out0;
wire  [14:0] v$_10659_out0;
wire  [14:0] v$_10660_out0;
wire  [14:0] v$_10661_out0;
wire  [14:0] v$_10662_out0;
wire  [14:0] v$_10663_out0;
wire  [14:0] v$_10664_out0;
wire  [14:0] v$_10665_out0;
wire  [14:0] v$_10666_out0;
wire  [14:0] v$_10667_out0;
wire  [14:0] v$_10668_out0;
wire  [14:0] v$_10669_out0;
wire  [14:0] v$_10670_out0;
wire  [14:0] v$_10671_out0;
wire  [14:0] v$_10672_out0;
wire  [14:0] v$_10673_out0;
wire  [14:0] v$_10674_out0;
wire  [14:0] v$_10675_out0;
wire  [14:0] v$_10676_out0;
wire  [14:0] v$_10677_out0;
wire  [14:0] v$_10678_out0;
wire  [14:0] v$_10679_out0;
wire  [14:0] v$_10680_out0;
wire  [14:0] v$_10910_out1;
wire  [14:0] v$_10911_out1;
wire  [14:0] v$_11231_out0;
wire  [14:0] v$_11232_out0;
wire  [14:0] v$_11294_out0;
wire  [14:0] v$_11295_out0;
wire  [14:0] v$_13709_out0;
wire  [14:0] v$_13710_out0;
wire  [14:0] v$_2223_out0;
wire  [14:0] v$_2224_out0;
wire  [14:0] v$_2889_out1;
wire  [14:0] v$_2890_out1;
wire  [14:0] v$_2984_out1;
wire  [14:0] v$_2985_out1;
wire  [14:0] v$_4831_out0;
wire  [14:0] v$_4832_out0;
wire  [14:0] v$_4856_out1;
wire  [14:0] v$_4857_out1;
wire  [15:0] v$16BIT$WORD$ANSWER_8821_out0;
wire  [15:0] v$16BIT$WORD$ANSWER_8822_out0;
wire  [15:0] v$A1_3174_out0;
wire  [15:0] v$A1_3175_out0;
wire  [15:0] v$A1_3855_out0;
wire  [15:0] v$A1_3856_out0;
wire  [15:0] v$A4_11227_out0;
wire  [15:0] v$A4_11228_out0;
wire  [15:0] v$A5_1901_out0;
wire  [15:0] v$A5_1902_out0;
wire  [15:0] v$A6_10463_out0;
wire  [15:0] v$A6_10464_out0;
wire  [15:0] v$A8_11155_out0;
wire  [15:0] v$A8_11156_out0;
wire  [15:0] v$ADDER$IN_8744_out0;
wire  [15:0] v$ADDER$IN_8745_out0;
wire  [15:0] v$ADDER$IN_8746_out0;
wire  [15:0] v$ADDER$IN_8747_out0;
wire  [15:0] v$ALUOUT_10528_out0;
wire  [15:0] v$ALUOUT_10529_out0;
wire  [15:0] v$ALUOUT_11053_out0;
wire  [15:0] v$ALUOUT_11054_out0;
wire  [15:0] v$ALUOUT_4494_out0;
wire  [15:0] v$ALUOUT_4495_out0;
wire  [15:0] v$ALUOUT_4607_out0;
wire  [15:0] v$ALUOUT_4608_out0;
wire  [15:0] v$ALUOUT_8856_out0;
wire  [15:0] v$ALUOUT_8857_out0;
wire  [15:0] v$ANDOUT_630_out0;
wire  [15:0] v$ANDOUT_631_out0;
wire  [15:0] v$ANDOUT_632_out0;
wire  [15:0] v$ANDOUT_633_out0;
wire  [15:0] v$A_10274_out0;
wire  [15:0] v$A_10275_out0;
wire  [15:0] v$A_10276_out0;
wire  [15:0] v$A_10277_out0;
wire  [15:0] v$A_11250_out0;
wire  [15:0] v$A_11251_out0;
wire  [15:0] v$A_11252_out0;
wire  [15:0] v$A_11253_out0;
wire  [15:0] v$B_3350_out0;
wire  [15:0] v$B_3352_out0;
wire  [15:0] v$C11_4539_out0;
wire  [15:0] v$C11_4540_out0;
wire  [15:0] v$C13_2185_out0;
wire  [15:0] v$C13_2186_out0;
wire  [15:0] v$C15_1730_out0;
wire  [15:0] v$C15_1731_out0;
wire  [15:0] v$C5_2688_out0;
wire  [15:0] v$C5_2689_out0;
wire  [15:0] v$C7_1865_out0;
wire  [15:0] v$C7_1866_out0;
wire  [15:0] v$CIN_2355_out0;
wire  [15:0] v$CIN_2357_out0;
wire  [15:0] v$CIN_2358_out0;
wire  [15:0] v$CIN_2359_out0;
wire  [15:0] v$CIN_2360_out0;
wire  [15:0] v$CIN_2361_out0;
wire  [15:0] v$CIN_2362_out0;
wire  [15:0] v$CIN_2363_out0;
wire  [15:0] v$CIN_2364_out0;
wire  [15:0] v$CIN_2365_out0;
wire  [15:0] v$CIN_2366_out0;
wire  [15:0] v$CIN_2367_out0;
wire  [15:0] v$CIN_2368_out0;
wire  [15:0] v$CIN_2369_out0;
wire  [15:0] v$CIN_2370_out0;
wire  [15:0] v$CIN_2372_out0;
wire  [15:0] v$CIN_2373_out0;
wire  [15:0] v$CIN_2374_out0;
wire  [15:0] v$CIN_2375_out0;
wire  [15:0] v$CIN_2376_out0;
wire  [15:0] v$CIN_2377_out0;
wire  [15:0] v$CIN_2378_out0;
wire  [15:0] v$CIN_2379_out0;
wire  [15:0] v$CIN_2380_out0;
wire  [15:0] v$CIN_2381_out0;
wire  [15:0] v$CIN_2382_out0;
wire  [15:0] v$CIN_2383_out0;
wire  [15:0] v$CIN_2384_out0;
wire  [15:0] v$COUT_10916_out0;
wire  [15:0] v$COUT_10917_out0;
wire  [15:0] v$COUT_10918_out0;
wire  [15:0] v$COUT_10919_out0;
wire  [15:0] v$COUT_10920_out0;
wire  [15:0] v$COUT_10921_out0;
wire  [15:0] v$COUT_10922_out0;
wire  [15:0] v$COUT_10923_out0;
wire  [15:0] v$COUT_10924_out0;
wire  [15:0] v$COUT_10925_out0;
wire  [15:0] v$COUT_10926_out0;
wire  [15:0] v$COUT_10927_out0;
wire  [15:0] v$COUT_10928_out0;
wire  [15:0] v$COUT_10929_out0;
wire  [15:0] v$COUT_10930_out0;
wire  [15:0] v$COUT_10931_out0;
wire  [15:0] v$COUT_10932_out0;
wire  [15:0] v$COUT_10933_out0;
wire  [15:0] v$COUT_10934_out0;
wire  [15:0] v$COUT_10935_out0;
wire  [15:0] v$COUT_10936_out0;
wire  [15:0] v$COUT_10937_out0;
wire  [15:0] v$COUT_10938_out0;
wire  [15:0] v$COUT_10939_out0;
wire  [15:0] v$COUT_10940_out0;
wire  [15:0] v$COUT_10941_out0;
wire  [15:0] v$COUT_10942_out0;
wire  [15:0] v$COUT_10943_out0;
wire  [15:0] v$COUT_10944_out0;
wire  [15:0] v$COUT_10945_out0;
wire  [15:0] v$DATA$IN_10552_out0;
wire  [15:0] v$DATA$IN_10553_out0;
wire  [15:0] v$DATA$OUT_1135_out0;
wire  [15:0] v$DATA$RAM$IN0_284_out0;
wire  [15:0] v$DATA$RAM$IN1_4779_out0;
wire  [15:0] v$DATA$RAM$IN_558_out0;
wire  [15:0] v$DATA$RAM$IN_559_out0;
wire  [15:0] v$DATA$to$transmit_4546_out0;
wire  [15:0] v$DATA0_13293_out0;
wire  [15:0] v$DATA0_4737_out0;
wire  [15:0] v$DATA1_1974_out0;
wire  [15:0] v$DATA1_603_out0;
wire  [15:0] v$DATA_10445_out0;
wire  [15:0] v$DATA_2469_out0;
wire  [15:0] v$DFQDF_3025_out0;
wire  [15:0] v$DFQDF_3026_out0;
wire  [15:0] v$DIN3_10310_out0;
wire  [15:0] v$DIN3_10311_out0;
wire  [15:0] v$DIN_2266_out0;
wire  [15:0] v$DIN_2267_out0;
wire  [15:0] v$DIN_9798_out0;
wire  [15:0] v$DIN_9799_out0;
wire  [15:0] v$DOUT1_1207_out0;
wire  [15:0] v$DOUT1_1208_out0;
wire  [15:0] v$DOUT2_1733_out0;
wire  [15:0] v$DOUT2_1734_out0;
wire  [15:0] v$FLOATING$REGISTER$IN_562_out0;
wire  [15:0] v$FLOATING$REGISTER$IN_563_out0;
wire  [15:0] v$IN_10403_out0;
wire  [15:0] v$IN_10404_out0;
wire  [15:0] v$IN_11258_out0;
wire  [15:0] v$IN_11259_out0;
wire  [15:0] v$IN_13306_out0;
wire  [15:0] v$IN_13307_out0;
wire  [15:0] v$IN_13548_out0;
wire  [15:0] v$IN_13549_out0;
wire  [15:0] v$IN_13788_out0;
wire  [15:0] v$IN_13789_out0;
wire  [15:0] v$IN_190_out0;
wire  [15:0] v$IN_191_out0;
wire  [15:0] v$IN_1964_out0;
wire  [15:0] v$IN_1965_out0;
wire  [15:0] v$IN_2350_out0;
wire  [15:0] v$IN_2351_out0;
wire  [15:0] v$IN_2664_out0;
wire  [15:0] v$IN_2665_out0;
wire  [15:0] v$IN_5796_out0;
wire  [15:0] v$IN_5797_out0;
wire  [15:0] v$IN_685_out0;
wire  [15:0] v$IN_686_out0;
wire  [15:0] v$IN_8838_out0;
wire  [15:0] v$IN_8839_out0;
wire  [15:0] v$IN_98_out0;
wire  [15:0] v$IN_99_out0;
wire  [15:0] v$IR_105_out0;
wire  [15:0] v$IR_106_out0;
wire  [15:0] v$IR_10816_out0;
wire  [15:0] v$IR_10817_out0;
wire  [15:0] v$IR_13480_out0;
wire  [15:0] v$IR_13481_out0;
wire  [15:0] v$IR_1871_out0;
wire  [15:0] v$IR_1872_out0;
wire  [15:0] v$IR_2826_out0;
wire  [15:0] v$IR_2827_out0;
wire  [15:0] v$IR_2901_out0;
wire  [15:0] v$IR_2902_out0;
wire  [15:0] v$IR_640_out0;
wire  [15:0] v$IR_641_out0;
wire  [15:0] v$IR_7112_out0;
wire  [15:0] v$IR_7113_out0;
wire  [15:0] v$IR_7706_out0;
wire  [15:0] v$IR_7707_out0;
wire  [15:0] v$KEXTEND_13329_out0;
wire  [15:0] v$KEXTEND_13330_out0;
wire  [15:0] v$LS$REGIN_3303_out0;
wire  [15:0] v$LS$REGIN_3304_out0;
wire  [15:0] v$M$REGIN_271_out0;
wire  [15:0] v$M$REGIN_272_out0;
wire  [15:0] v$MEM$RAM_434_out0;
wire  [15:0] v$MEM$RAM_435_out0;
wire  [15:0] v$MULTI$OUT_13607_out0;
wire  [15:0] v$MULTI$OUT_13608_out0;
wire  [15:0] v$MULTI$OUT_1669_out0;
wire  [15:0] v$MULTI$OUT_1670_out0;
wire  [15:0] v$MULTI$REGIN_2870_out0;
wire  [15:0] v$MULTI$REGIN_2871_out0;
wire  [15:0] v$MUX11_13745_out0;
wire  [15:0] v$MUX11_13746_out0;
wire  [15:0] v$MUX12_1714_out0;
wire  [15:0] v$MUX12_1715_out0;
wire  [15:0] v$MUX1_10443_out0;
wire  [15:0] v$MUX1_10444_out0;
wire  [15:0] v$MUX1_11141_out0;
wire  [15:0] v$MUX1_11142_out0;
wire  [15:0] v$MUX1_1735_out0;
wire  [15:0] v$MUX1_1736_out0;
wire  [15:0] v$MUX1_1883_out0;
wire  [15:0] v$MUX1_1884_out0;
wire  [15:0] v$MUX1_2532_out0;
wire  [15:0] v$MUX1_2533_out0;
wire  [15:0] v$MUX1_2717_out0;
wire  [15:0] v$MUX1_2718_out0;
wire  [15:0] v$MUX1_31_out0;
wire  [15:0] v$MUX1_32_out0;
wire  [15:0] v$MUX1_4844_out0;
wire  [15:0] v$MUX1_4845_out0;
wire  [15:0] v$MUX1_6_out0;
wire  [15:0] v$MUX1_7_out0;
wire  [15:0] v$MUX1_8813_out0;
wire  [15:0] v$MUX1_8814_out0;
wire  [15:0] v$MUX2_10841_out0;
wire  [15:0] v$MUX2_10842_out0;
wire  [15:0] v$MUX2_1181_out0;
wire  [15:0] v$MUX2_1182_out0;
wire  [15:0] v$MUX2_1199_out0;
wire  [15:0] v$MUX2_1200_out0;
wire  [15:0] v$MUX2_13319_out0;
wire  [15:0] v$MUX2_13320_out0;
wire  [15:0] v$MUX2_2337_out0;
wire  [15:0] v$MUX2_2338_out0;
wire  [15:0] v$MUX2_3202_out0;
wire  [15:0] v$MUX2_3203_out0;
wire  [15:0] v$MUX2_3255_out0;
wire  [15:0] v$MUX2_3256_out0;
wire  [15:0] v$MUX2_4612_out0;
wire  [15:0] v$MUX2_4613_out0;
wire  [15:0] v$MUX3_10787_out0;
wire  [15:0] v$MUX3_13335_out0;
wire  [15:0] v$MUX3_13336_out0;
wire  [15:0] v$MUX3_2058_out0;
wire  [15:0] v$MUX3_2059_out0;
wire  [15:0] v$MUX3_3041_out0;
wire  [15:0] v$MUX3_3042_out0;
wire  [15:0] v$MUX3_3133_out0;
wire  [15:0] v$MUX3_3134_out0;
wire  [15:0] v$MUX3_313_out0;
wire  [15:0] v$MUX3_314_out0;
wire  [15:0] v$MUX3_6864_out0;
wire  [15:0] v$MUX3_6865_out0;
wire  [15:0] v$MUX3_7075_out0;
wire  [15:0] v$MUX3_7076_out0;
wire  [15:0] v$MUX3_8669_out0;
wire  [15:0] v$MUX3_8670_out0;
wire  [15:0] v$MUX4_10524_out0;
wire  [15:0] v$MUX4_10525_out0;
wire  [15:0] v$MUX4_10_out0;
wire  [15:0] v$MUX4_11_out0;
wire  [15:0] v$MUX4_13498_out0;
wire  [15:0] v$MUX4_13499_out0;
wire  [15:0] v$MUX4_1698_out0;
wire  [15:0] v$MUX4_2229_out0;
wire  [15:0] v$MUX4_2230_out0;
wire  [15:0] v$MUX4_376_out0;
wire  [15:0] v$MUX4_377_out0;
wire  [15:0] v$MUX4_4579_out0;
wire  [15:0] v$MUX4_4580_out0;
wire  [15:0] v$MUX4_7023_out0;
wire  [15:0] v$MUX4_7024_out0;
wire  [15:0] v$MUX5_10605_out0;
wire  [15:0] v$MUX5_10606_out0;
wire  [15:0] v$MUX5_1185_out0;
wire  [15:0] v$MUX5_1186_out0;
wire  [15:0] v$MUX5_2595_out0;
wire  [15:0] v$MUX5_2596_out0;
wire  [15:0] v$MUX5_2606_out0;
wire  [15:0] v$MUX5_2607_out0;
wire  [15:0] v$MUX5_3305_out0;
wire  [15:0] v$MUX5_3306_out0;
wire  [15:0] v$MUX5_7017_out0;
wire  [15:0] v$MUX5_7018_out0;
wire  [15:0] v$MUX5_8840_out0;
wire  [15:0] v$MUX5_8841_out0;
wire  [15:0] v$MUX6_2341_out0;
wire  [15:0] v$MUX6_2342_out0;
wire  [15:0] v$MUX7_1165_out0;
wire  [15:0] v$MUX7_1166_out0;
wire  [15:0] v$MUX8_1907_out0;
wire  [15:0] v$MUX8_1908_out0;
wire  [15:0] v$OP1_2060_out0;
wire  [15:0] v$OP1_2061_out0;
wire  [15:0] v$OP1_2979_out0;
wire  [15:0] v$OP1_2980_out0;
wire  [15:0] v$OP1_3899_out0;
wire  [15:0] v$OP1_3900_out0;
wire  [15:0] v$OP2_10751_out0;
wire  [15:0] v$OP2_10752_out0;
wire  [15:0] v$OP2_11153_out0;
wire  [15:0] v$OP2_11154_out0;
wire  [15:0] v$OP2_2322_out0;
wire  [15:0] v$OP2_2323_out0;
wire  [15:0] v$OP2_2862_out0;
wire  [15:0] v$OP2_2863_out0;
wire  [15:0] v$OP2_3940_out0;
wire  [15:0] v$OP2_3941_out0;
wire  [15:0] v$OUT_10264_out0;
wire  [15:0] v$OUT_10265_out0;
wire  [15:0] v$OUT_11234_out0;
wire  [15:0] v$OUT_11235_out0;
wire  [15:0] v$OUT_1136_out0;
wire  [15:0] v$OUT_1137_out0;
wire  [15:0] v$OUT_12236_out0;
wire  [15:0] v$OUT_12237_out0;
wire  [15:0] v$OUT_2352_out0;
wire  [15:0] v$OUT_2353_out0;
wire  [15:0] v$OUT_2857_out0;
wire  [15:0] v$OUT_2858_out0;
wire  [15:0] v$OUT_460_out0;
wire  [15:0] v$OUT_461_out0;
wire  [15:0] v$OUT_7708_out0;
wire  [15:0] v$OUT_7709_out0;
wire  [15:0] v$OUT_7710_out0;
wire  [15:0] v$OUT_7711_out0;
wire  [15:0] v$OUT_8852_out0;
wire  [15:0] v$OUT_8853_out0;
wire  [15:0] v$R0TEST_3184_out0;
wire  [15:0] v$R0TEST_3185_out0;
wire  [15:0] v$R0TEST_7005_out0;
wire  [15:0] v$R0TEST_7006_out0;
wire  [15:0] v$R0_13295_out0;
wire  [15:0] v$R0_13296_out0;
wire  [15:0] v$R0_1688_out0;
wire  [15:0] v$R0_1689_out0;
wire  [15:0] v$R0_2537_out0;
wire  [15:0] v$R0_2538_out0;
wire  [15:0] v$R0_2850_out0;
wire  [15:0] v$R0_2851_out0;
wire  [15:0] v$R1TEST_10485_out0;
wire  [15:0] v$R1TEST_10486_out0;
wire  [15:0] v$R1TEST_10498_out0;
wire  [15:0] v$R1TEST_10499_out0;
wire  [15:0] v$R1_2056_out0;
wire  [15:0] v$R1_2057_out0;
wire  [15:0] v$R1_2630_out0;
wire  [15:0] v$R1_2631_out0;
wire  [15:0] v$R1_2723_out0;
wire  [15:0] v$R1_2724_out0;
wire  [15:0] v$R1_8761_out0;
wire  [15:0] v$R1_8762_out0;
wire  [15:0] v$R2TEST_10708_out0;
wire  [15:0] v$R2TEST_10709_out0;
wire  [15:0] v$R2TEST_10987_out0;
wire  [15:0] v$R2TEST_10988_out0;
wire  [15:0] v$R2_10556_out0;
wire  [15:0] v$R2_10557_out0;
wire  [15:0] v$R2_10904_out0;
wire  [15:0] v$R2_10905_out0;
wire  [15:0] v$R2_1726_out0;
wire  [15:0] v$R2_1727_out0;
wire  [15:0] v$R2_3043_out0;
wire  [15:0] v$R2_3044_out0;
wire  [15:0] v$R3TEST_117_out0;
wire  [15:0] v$R3TEST_118_out0;
wire  [15:0] v$R3TEST_2872_out0;
wire  [15:0] v$R3TEST_2873_out0;
wire  [15:0] v$R3_27_out0;
wire  [15:0] v$R3_28_out0;
wire  [15:0] v$R3_33_out0;
wire  [15:0] v$R3_34_out0;
wire  [15:0] v$R3_4652_out0;
wire  [15:0] v$R3_4653_out0;
wire  [15:0] v$R3_74_out0;
wire  [15:0] v$R3_75_out0;
wire  [15:0] v$RAM$IN_233_out0;
wire  [15:0] v$RAM$IN_234_out0;
wire  [15:0] v$RAM$OUT0_8764_out0;
wire  [15:0] v$RAM$OUT1_2385_out0;
wire  [15:0] v$RAM$OUT_10335_out0;
wire  [15:0] v$RAM$OUT_10336_out0;
wire  [15:0] v$RAM$OUT_11214_out0;
wire  [15:0] v$RAM$OUT_11215_out0;
wire  [15:0] v$RAM$OUT_1751_out0;
wire  [15:0] v$RAM$OUT_1752_out0;
wire  [15:0] v$RAM$OUT_2104_out0;
wire  [15:0] v$RAM$OUT_2105_out0;
wire  [15:0] v$RAM$OUT_2628_out0;
wire  [15:0] v$RAM$OUT_2629_out0;
wire  [15:0] v$RAM$OUT_3033_out0;
wire  [15:0] v$RAM$OUT_3034_out0;
wire  [15:0] v$RAM0_1680_out0;
wire  [15:0] v$RAM1_13398_out0;
wire  [15:0] v$RAMDOUT_23_out0;
wire  [15:0] v$RAMDOUT_2414_out0;
wire  [15:0] v$RAMDOUT_2415_out0;
wire  [15:0] v$RAMDOUT_24_out0;
wire  [15:0] v$RAMDOUT_3031_out0;
wire  [15:0] v$RAMDOUT_3032_out0;
wire  [15:0] v$RD$FLOATING_2823_out0;
wire  [15:0] v$RD$FLOATING_2824_out0;
wire  [15:0] v$RD$MULTI_45_out0;
wire  [15:0] v$RD$MULTI_46_out0;
wire  [15:0] v$RD$STATUS_10500_out0;
wire  [15:0] v$RDOUT_2787_out0;
wire  [15:0] v$RDOUT_2788_out0;
wire  [15:0] v$RD_3891_out0;
wire  [15:0] v$RD_3892_out0;
wire  [15:0] v$RD_4839_out0;
wire  [15:0] v$RD_4840_out0;
wire  [15:0] v$RD_501_out0;
wire  [15:0] v$RD_502_out0;
wire  [15:0] v$RD_613_out0;
wire  [15:0] v$RD_614_out0;
wire  [15:0] v$REGDIN_11041_out0;
wire  [15:0] v$REGDIN_11042_out0;
wire  [15:0] v$REGISTE$IN_4490_out0;
wire  [15:0] v$REGISTE$IN_4491_out0;
wire  [15:0] v$REGISTER$INPUT_13270_out0;
wire  [15:0] v$REGISTER$INPUT_13271_out0;
wire  [15:0] v$REGISTER$INPUT_13621_out0;
wire  [15:0] v$REGISTER$INPUT_13622_out0;
wire  [15:0] v$REGISTER$OUTPUT2_2398_out0;
wire  [15:0] v$REGISTER$OUTPUT_3268_out0;
wire  [15:0] v$REGISTER$OUT_10268_out0;
wire  [15:0] v$REGISTER$OUT_10269_out0;
wire  [15:0] v$RM$MULTI_210_out0;
wire  [15:0] v$RM$MULTI_211_out0;
wire  [15:0] v$RM$MULTI_648_out0;
wire  [15:0] v$RM$MULTI_649_out0;
wire  [15:0] v$RMN_13437_out0;
wire  [15:0] v$RMN_13438_out0;
wire  [15:0] v$RM_11063_out0;
wire  [15:0] v$RM_11064_out0;
wire  [15:0] v$RM_11065_out0;
wire  [15:0] v$RM_11066_out0;
wire  [15:0] v$RM_11067_out0;
wire  [15:0] v$RM_11068_out0;
wire  [15:0] v$RM_11069_out0;
wire  [15:0] v$RM_11070_out0;
wire  [15:0] v$RM_11071_out0;
wire  [15:0] v$RM_11072_out0;
wire  [15:0] v$RM_11073_out0;
wire  [15:0] v$RM_11074_out0;
wire  [15:0] v$RM_11075_out0;
wire  [15:0] v$RM_11076_out0;
wire  [15:0] v$RM_11077_out0;
wire  [15:0] v$RM_11078_out0;
wire  [15:0] v$RM_11079_out0;
wire  [15:0] v$RM_11080_out0;
wire  [15:0] v$RM_11081_out0;
wire  [15:0] v$RM_11082_out0;
wire  [15:0] v$RM_11083_out0;
wire  [15:0] v$RM_11084_out0;
wire  [15:0] v$RM_11085_out0;
wire  [15:0] v$RM_11086_out0;
wire  [15:0] v$RM_11087_out0;
wire  [15:0] v$RM_11088_out0;
wire  [15:0] v$RM_11089_out0;
wire  [15:0] v$RM_11090_out0;
wire  [15:0] v$RM_11091_out0;
wire  [15:0] v$RM_11092_out0;
wire  [15:0] v$RM_11167_out0;
wire  [15:0] v$RM_11168_out0;
wire  [15:0] v$RM_13508_out0;
wire  [15:0] v$RM_13509_out0;
wire  [15:0] v$RM_13597_out0;
wire  [15:0] v$RM_13598_out0;
wire  [15:0] v$RM_13750_out0;
wire  [15:0] v$RM_13751_out0;
wire  [15:0] v$RM_2432_out0;
wire  [15:0] v$RM_2433_out0;
wire  [15:0] v$RM_2912_out0;
wire  [15:0] v$RM_2913_out0;
wire  [15:0] v$RM_3272_out0;
wire  [15:0] v$RM_3273_out0;
wire  [15:0] v$RM_4537_out0;
wire  [15:0] v$RM_4538_out0;
wire  [15:0] v$RM_8731_out0;
wire  [15:0] v$RM_8732_out0;
wire  [15:0] v$STATUS$REGISTER_10359_out0;
wire  [15:0] v$STATUS$REGISTER_13778_out0;
wire  [15:0] v$STATUS$REGISTER_185_out0;
wire  [15:0] v$STATUS$REGISTER_2866_out0;
wire  [15:0] v$STATUS$REGISTER_2867_out0;
wire  [15:0] v$STATUS$REGISTER_5858_out0;
wire  [15:0] v$STATUS$REGISTER_5859_out0;
wire  [15:0] v$SUM1_13213_out0;
wire  [15:0] v$SUM1_13214_out0;
wire  [15:0] v$XOR1_11246_out0;
wire  [15:0] v$XOR1_11247_out0;
wire  [15:0] v$XOR2_4486_out0;
wire  [15:0] v$XOR2_4487_out0;
wire  [15:0] v$XOR3_13599_out0;
wire  [15:0] v$XOR3_13600_out0;
wire  [15:0] v$_10333_out0;
wire  [15:0] v$_10334_out0;
wire  [15:0] v$_10449_out0;
wire  [15:0] v$_10450_out0;
wire  [15:0] v$_10504_out0;
wire  [15:0] v$_10505_out0;
wire  [15:0] v$_10532_out0;
wire  [15:0] v$_10814_out0;
wire  [15:0] v$_10815_out0;
wire  [15:0] v$_10946_out0;
wire  [15:0] v$_10947_out0;
wire  [15:0] v$_10948_out0;
wire  [15:0] v$_10949_out0;
wire  [15:0] v$_10950_out0;
wire  [15:0] v$_10951_out0;
wire  [15:0] v$_10952_out0;
wire  [15:0] v$_10953_out0;
wire  [15:0] v$_10954_out0;
wire  [15:0] v$_10955_out0;
wire  [15:0] v$_10956_out0;
wire  [15:0] v$_10957_out0;
wire  [15:0] v$_10958_out0;
wire  [15:0] v$_10959_out0;
wire  [15:0] v$_10960_out0;
wire  [15:0] v$_10961_out0;
wire  [15:0] v$_10962_out0;
wire  [15:0] v$_10963_out0;
wire  [15:0] v$_10964_out0;
wire  [15:0] v$_10965_out0;
wire  [15:0] v$_10966_out0;
wire  [15:0] v$_10967_out0;
wire  [15:0] v$_10968_out0;
wire  [15:0] v$_10969_out0;
wire  [15:0] v$_10970_out0;
wire  [15:0] v$_10971_out0;
wire  [15:0] v$_10972_out0;
wire  [15:0] v$_10973_out0;
wire  [15:0] v$_10974_out0;
wire  [15:0] v$_10975_out0;
wire  [15:0] v$_11229_out0;
wire  [15:0] v$_11230_out0;
wire  [15:0] v$_1172_out0;
wire  [15:0] v$_1173_out0;
wire  [15:0] v$_1209_out0;
wire  [15:0] v$_1210_out0;
wire  [15:0] v$_1211_out0;
wire  [15:0] v$_1212_out0;
wire  [15:0] v$_1213_out0;
wire  [15:0] v$_1214_out0;
wire  [15:0] v$_124_out0;
wire  [15:0] v$_125_out0;
wire  [15:0] v$_13275_out0;
wire  [15:0] v$_13276_out0;
wire  [15:0] v$_13482_out0;
wire  [15:0] v$_13483_out0;
wire  [15:0] v$_167_out0;
wire  [15:0] v$_168_out0;
wire  [15:0] v$_1867_out0;
wire  [15:0] v$_1868_out0;
wire  [15:0] v$_1869_out0;
wire  [15:0] v$_1870_out0;
wire  [15:0] v$_2678_out0;
wire  [15:0] v$_2679_out0;
wire  [15:0] v$_2791_out0;
wire  [15:0] v$_2792_out0;
wire  [15:0] v$_3178_out0;
wire  [15:0] v$_3179_out0;
wire  [15:0] v$_333_out0;
wire  [15:0] v$_334_out0;
wire  [15:0] v$_403_out0;
wire  [15:0] v$_404_out0;
wire  [15:0] v$_4660_out0;
wire  [15:0] v$_4661_out0;
wire  [15:0] v$_4709_out0;
wire  [15:0] v$_4710_out0;
wire  [15:0] v$_6870_out0;
wire  [15:0] v$_6871_out0;
wire  [15:0] v$_7081_out0;
wire  [15:0] v$_7082_out0;
wire  [15:0] v$_7120_out0;
wire  [15:0] v$_7121_out0;
wire  [15:0] v$_7124_out0;
wire  [15:0] v$_7125_out0;
wire  [15:0] v$_7179_out0;
wire  [15:0] v$_7180_out0;
wire  [15:0] v$_7638_out0;
wire  [15:0] v$_7639_out0;
wire  [15:0] v$_7640_out0;
wire  [15:0] v$_7641_out0;
wire  [15:0] v$_8697_out0;
wire  [15:0] v$_8698_out0;
wire  [15:0] v$_9791_out0;
wire  [15:0] v$_9792_out0;
wire  [15:0] v$data$ram_1818_out0;
wire  [1:0] v$4BITCOUNTER_317_out0;
wire  [1:0] v$4BITCOUNTER_318_out0;
wire  [1:0] v$4BITCOUNTER_319_out0;
wire  [1:0] v$4BITCOUNTER_320_out0;
wire  [1:0] v$AD1_13774_out0;
wire  [1:0] v$AD1_13775_out0;
wire  [1:0] v$AD2_10699_out0;
wire  [1:0] v$AD2_10700_out0;
wire  [1:0] v$AD3_10482_out0;
wire  [1:0] v$AD3_10483_out0;
wire  [1:0] v$AD3_13272_out0;
wire  [1:0] v$AD3_13273_out0;
wire  [1:0] v$AD3_8671_out0;
wire  [1:0] v$AD3_8672_out0;
wire  [1:0] v$C1_11292_out0;
wire  [1:0] v$C1_11293_out0;
wire  [1:0] v$C1_3205_out0;
wire  [1:0] v$C1_3206_out0;
wire  [1:0] v$C1_6793_out0;
wire  [1:0] v$C1_6794_out0;
wire  [1:0] v$C5_10356_out0;
wire  [1:0] v$D_2108_out0;
wire  [1:0] v$D_2109_out0;
wire  [1:0] v$D_623_out0;
wire  [1:0] v$D_624_out0;
wire  [1:0] v$D_8752_out0;
wire  [1:0] v$D_8753_out0;
wire  [1:0] v$MUX1_11061_out0;
wire  [1:0] v$MUX1_534_out0;
wire  [1:0] v$MUX1_535_out0;
wire  [1:0] v$MUX2_1145_out0;
wire  [1:0] v$MUX2_1146_out0;
wire  [1:0] v$M_4701_out0;
wire  [1:0] v$M_4702_out0;
wire  [1:0] v$M_7177_out0;
wire  [1:0] v$M_7178_out0;
wire  [1:0] v$NOTUSED_2589_out0;
wire  [1:0] v$NOTUSED_2590_out0;
wire  [1:0] v$NOTUSED_445_out0;
wire  [1:0] v$NOTUSED_446_out0;
wire  [1:0] v$NOTUSED_447_out0;
wire  [1:0] v$NOTUSED_448_out0;
wire  [1:0] v$Q_10618_out0;
wire  [1:0] v$Q_1153_out0;
wire  [1:0] v$Q_1154_out0;
wire  [1:0] v$Q_13510_out0;
wire  [1:0] v$RD_10522_out0;
wire  [1:0] v$RD_10523_out0;
wire  [1:0] v$ROR_66_out0;
wire  [1:0] v$ROR_67_out0;
wire  [1:0] v$SHIFT_10615_out0;
wire  [1:0] v$SHIFT_10616_out0;
wire  [1:0] v$SHIFT_8661_out0;
wire  [1:0] v$SHIFT_8662_out0;
wire  [1:0] v$SR_10607_out0;
wire  [1:0] v$SR_10608_out0;
wire  [1:0] v$SR_1956_out0;
wire  [1:0] v$SR_1957_out0;
wire  [1:0] v$SR_371_out0;
wire  [1:0] v$SR_372_out0;
wire  [1:0] v$SR_542_out0;
wire  [1:0] v$SR_543_out0;
wire  [1:0] v$UNUSED_11244_out0;
wire  [1:0] v$UNUSED_11245_out0;
wire  [1:0] v$_10287_out0;
wire  [1:0] v$_10288_out0;
wire  [1:0] v$_10289_out0;
wire  [1:0] v$_10290_out0;
wire  [1:0] v$_10791_out0;
wire  [1:0] v$_10792_out0;
wire  [1:0] v$_11049_out1;
wire  [1:0] v$_11050_out1;
wire  [1:0] v$_11057_out0;
wire  [1:0] v$_11058_out0;
wire  [1:0] v$_11163_out0;
wire  [1:0] v$_11164_out0;
wire  [1:0] v$_1140_out0;
wire  [1:0] v$_1141_out0;
wire  [1:0] v$_13261_out0;
wire  [1:0] v$_13262_out0;
wire  [1:0] v$_13263_out0;
wire  [1:0] v$_13264_out0;
wire  [1:0] v$_13550_out0;
wire  [1:0] v$_13551_out0;
wire  [1:0] v$_13770_out0;
wire  [1:0] v$_13771_out0;
wire  [1:0] v$_13772_out0;
wire  [1:0] v$_13773_out0;
wire  [1:0] v$_1707_out0;
wire  [1:0] v$_1708_out0;
wire  [1:0] v$_1951_out0;
wire  [1:0] v$_1952_out0;
wire  [1:0] v$_1953_out0;
wire  [1:0] v$_1954_out0;
wire  [1:0] v$_2599_out0;
wire  [1:0] v$_2600_out0;
wire  [1:0] v$_2887_out0;
wire  [1:0] v$_2888_out0;
wire  [1:0] v$_2945_out0;
wire  [1:0] v$_2946_out0;
wire  [1:0] v$_2947_out0;
wire  [1:0] v$_2948_out0;
wire  [1:0] v$_3215_out0;
wire  [1:0] v$_3216_out0;
wire  [1:0] v$_3217_out0;
wire  [1:0] v$_3218_out0;
wire  [1:0] v$_3223_out0;
wire  [1:0] v$_3224_out0;
wire  [1:0] v$_3278_out0;
wire  [1:0] v$_3279_out0;
wire  [1:0] v$_3280_out0;
wire  [1:0] v$_3281_out0;
wire  [1:0] v$_386_out0;
wire  [1:0] v$_387_out0;
wire  [1:0] v$_388_out0;
wire  [1:0] v$_389_out0;
wire  [1:0] v$_399_out0;
wire  [1:0] v$_400_out0;
wire  [1:0] v$_401_out0;
wire  [1:0] v$_402_out0;
wire  [1:0] v$_4483_out0;
wire  [1:0] v$_4484_out0;
wire  [1:0] v$_4547_out0;
wire  [1:0] v$_4782_out0;
wire  [1:0] v$_4783_out0;
wire  [1:0] v$_4784_out0;
wire  [1:0] v$_4785_out0;
wire  [1:0] v$_4786_out0;
wire  [1:0] v$_4787_out0;
wire  [1:0] v$_4788_out0;
wire  [1:0] v$_4789_out0;
wire  [1:0] v$_4790_out0;
wire  [1:0] v$_4791_out0;
wire  [1:0] v$_4792_out0;
wire  [1:0] v$_4793_out0;
wire  [1:0] v$_4794_out0;
wire  [1:0] v$_4795_out0;
wire  [1:0] v$_4796_out0;
wire  [1:0] v$_4797_out0;
wire  [1:0] v$_4798_out0;
wire  [1:0] v$_4799_out0;
wire  [1:0] v$_4800_out0;
wire  [1:0] v$_4801_out0;
wire  [1:0] v$_4802_out0;
wire  [1:0] v$_4803_out0;
wire  [1:0] v$_4804_out0;
wire  [1:0] v$_4805_out0;
wire  [1:0] v$_4806_out0;
wire  [1:0] v$_4807_out0;
wire  [1:0] v$_4808_out0;
wire  [1:0] v$_4809_out0;
wire  [1:0] v$_4810_out0;
wire  [1:0] v$_4811_out0;
wire  [1:0] v$_4816_out0;
wire  [1:0] v$_4817_out0;
wire  [1:0] v$_533_out0;
wire  [1:0] v$_627_out0;
wire  [1:0] v$_628_out0;
wire  [1:0] v$_7135_out0;
wire  [1:0] v$_7136_out0;
wire  [1:0] v$_7137_out0;
wire  [1:0] v$_7138_out0;
wire  [1:0] v$_7183_out0;
wire  [1:0] v$_7184_out0;
wire  [1:0] v$_7185_out0;
wire  [1:0] v$_7186_out0;
wire  [2:0] v$C1_2716_out0;
wire  [2:0] v$C2_11233_out0;
wire  [2:0] v$C3_10853_out0;
wire  [2:0] v$C4_1201_out0;
wire  [2:0] v$OP_11223_out0;
wire  [2:0] v$OP_11224_out0;
wire  [2:0] v$OP_621_out0;
wire  [2:0] v$OP_622_out0;
wire  [2:0] v$_13253_out0;
wire  [2:0] v$_13254_out0;
wire  [2:0] v$_1716_out0;
wire  [2:0] v$_1717_out0;
wire  [2:0] v$_2386_out0;
wire  [2:0] v$_2387_out0;
wire  [2:0] v$_2552_out0;
wire  [2:0] v$_2553_out0;
wire  [2:0] v$_2554_out0;
wire  [2:0] v$_2555_out0;
wire  [2:0] v$_2556_out0;
wire  [2:0] v$_2557_out0;
wire  [2:0] v$_2558_out0;
wire  [2:0] v$_2559_out0;
wire  [2:0] v$_2560_out0;
wire  [2:0] v$_2561_out0;
wire  [2:0] v$_2562_out0;
wire  [2:0] v$_2563_out0;
wire  [2:0] v$_2564_out0;
wire  [2:0] v$_2565_out0;
wire  [2:0] v$_2566_out0;
wire  [2:0] v$_2567_out0;
wire  [2:0] v$_2568_out0;
wire  [2:0] v$_2569_out0;
wire  [2:0] v$_2570_out0;
wire  [2:0] v$_2571_out0;
wire  [2:0] v$_2572_out0;
wire  [2:0] v$_2573_out0;
wire  [2:0] v$_2574_out0;
wire  [2:0] v$_2575_out0;
wire  [2:0] v$_2576_out0;
wire  [2:0] v$_2577_out0;
wire  [2:0] v$_2578_out0;
wire  [2:0] v$_2579_out0;
wire  [2:0] v$_2580_out0;
wire  [2:0] v$_2581_out0;
wire  [2:0] v$_2680_out1;
wire  [2:0] v$_2681_out1;
wire  [2:0] v$_2960_out0;
wire  [2:0] v$_2961_out0;
wire  [2:0] v$_2962_out0;
wire  [2:0] v$_2963_out0;
wire  [2:0] v$_4_out0;
wire  [2:0] v$_5_out0;
wire  [2:0] v$_9804_out0;
wire  [2:0] v$_9805_out0;
wire  [2:0] v$_9806_out0;
wire  [2:0] v$_9807_out0;
wire  [31:0] v$32BIT$MULTI_1183_out0;
wire  [31:0] v$32BIT$MULTI_1184_out0;
wire  [31:0] v$32BITPRODUCT_12249_out0;
wire  [31:0] v$32BITPRODUCT_12250_out0;
wire  [31:0] v$32BITPRODUCT_82_out0;
wire  [31:0] v$32BITPRODUCT_83_out0;
wire  [31:0] v$FLOATING$MULTI_7697_out0;
wire  [31:0] v$FLOATING$MULTI_7698_out0;
wire  [31:0] v$_212_out0;
wire  [31:0] v$_213_out0;
wire  [3:0] v$8BITCOUNTER_13281_out0;
wire  [3:0] v$8BITCOUNTER_13282_out0;
wire  [3:0] v$8BITCOUNTER_13283_out0;
wire  [3:0] v$8BITCOUNTER_13284_out0;
wire  [3:0] v$BIN_5853_out0;
wire  [3:0] v$BIN_5854_out0;
wire  [3:0] v$B_10793_out0;
wire  [3:0] v$B_10794_out0;
wire  [3:0] v$B_1155_out0;
wire  [3:0] v$B_1156_out0;
wire  [3:0] v$B_273_out0;
wire  [3:0] v$B_274_out0;
wire  [3:0] v$C1_10305_out0;
wire  [3:0] v$C1_10306_out0;
wire  [3:0] v$C1_2005_out0;
wire  [3:0] v$C1_2006_out0;
wire  [3:0] v$C1_6919_out0;
wire  [3:0] v$C1_6920_out0;
wire  [3:0] v$MUX1_2409_out0;
wire  [3:0] v$MUX1_2410_out0;
wire  [3:0] v$NOTUSED1_1897_out0;
wire  [3:0] v$NOTUSED1_1898_out0;
wire  [3:0] v$NOTUSED_10540_out0;
wire  [3:0] v$NOTUSED_10541_out0;
wire  [3:0] v$NOTUSED_13265_out0;
wire  [3:0] v$NOTUSED_13266_out0;
wire  [3:0] v$NOTUSED_9800_out0;
wire  [3:0] v$NOTUSED_9801_out0;
wire  [3:0] v$NOTUSE_2399_out0;
wire  [3:0] v$NOTUSE_2400_out0;
wire  [3:0] v$N_7642_out0;
wire  [3:0] v$N_7643_out0;
wire  [3:0] v$RAM$ADD$BYTE0_13382_out0;
wire  [3:0] v$RAM$ADD$BYTE0_13383_out0;
wire  [3:0] v$SEL1_5798_out0;
wire  [3:0] v$SEL1_5799_out0;
wire  [3:0] v$UNUSED_13431_out0;
wire  [3:0] v$UNUSED_13432_out0;
wire  [3:0] v$_10372_out0;
wire  [3:0] v$_10373_out0;
wire  [3:0] v$_10374_out0;
wire  [3:0] v$_10375_out0;
wire  [3:0] v$_113_out0;
wire  [3:0] v$_1140_out1;
wire  [3:0] v$_1141_out1;
wire  [3:0] v$_114_out0;
wire  [3:0] v$_115_out0;
wire  [3:0] v$_116_out0;
wire  [3:0] v$_13291_out0;
wire  [3:0] v$_13292_out0;
wire  [3:0] v$_13317_out0;
wire  [3:0] v$_13317_out1;
wire  [3:0] v$_13318_out0;
wire  [3:0] v$_13318_out1;
wire  [3:0] v$_13337_out0;
wire  [3:0] v$_1673_out0;
wire  [3:0] v$_1813_out0;
wire  [3:0] v$_2146_out0;
wire  [3:0] v$_2147_out0;
wire  [3:0] v$_224_out1;
wire  [3:0] v$_225_out1;
wire  [3:0] v$_2345_out0;
wire  [3:0] v$_2346_out0;
wire  [3:0] v$_2347_out0;
wire  [3:0] v$_2348_out0;
wire  [3:0] v$_2411_out1;
wire  [3:0] v$_2412_out1;
wire  [3:0] v$_2437_out0;
wire  [3:0] v$_2438_out0;
wire  [3:0] v$_2536_out0;
wire  [3:0] v$_2773_out0;
wire  [3:0] v$_2774_out0;
wire  [3:0] v$_2775_out0;
wire  [3:0] v$_2776_out0;
wire  [3:0] v$_2968_out0;
wire  [3:0] v$_2969_out0;
wire  [3:0] v$_3035_out1;
wire  [3:0] v$_3036_out1;
wire  [3:0] v$_3942_out0;
wire  [3:0] v$_3943_out0;
wire  [3:0] v$_4488_out0;
wire  [3:0] v$_4489_out0;
wire  [3:0] v$_449_out0;
wire  [3:0] v$_450_out0;
wire  [3:0] v$_451_out0;
wire  [3:0] v$_4529_out0;
wire  [3:0] v$_452_out0;
wire  [3:0] v$_4530_out0;
wire  [3:0] v$_4585_out0;
wire  [3:0] v$_4586_out0;
wire  [3:0] v$_4703_out0;
wire  [3:0] v$_4704_out0;
wire  [3:0] v$_5846_out1;
wire  [3:0] v$_5847_out1;
wire  [3:0] v$_7032_out0;
wire  [3:0] v$_7033_out0;
wire  [3:0] v$_7034_out0;
wire  [3:0] v$_7035_out0;
wire  [3:0] v$_7036_out0;
wire  [3:0] v$_7037_out0;
wire  [3:0] v$_7038_out0;
wire  [3:0] v$_7039_out0;
wire  [3:0] v$_7040_out0;
wire  [3:0] v$_7041_out0;
wire  [3:0] v$_7042_out0;
wire  [3:0] v$_7043_out0;
wire  [3:0] v$_7044_out0;
wire  [3:0] v$_7045_out0;
wire  [3:0] v$_7046_out0;
wire  [3:0] v$_7047_out0;
wire  [3:0] v$_7048_out0;
wire  [3:0] v$_7049_out0;
wire  [3:0] v$_7050_out0;
wire  [3:0] v$_7051_out0;
wire  [3:0] v$_7052_out0;
wire  [3:0] v$_7053_out0;
wire  [3:0] v$_7054_out0;
wire  [3:0] v$_7055_out0;
wire  [3:0] v$_7056_out0;
wire  [3:0] v$_7057_out0;
wire  [3:0] v$_7058_out0;
wire  [3:0] v$_7059_out0;
wire  [3:0] v$_7060_out0;
wire  [3:0] v$_7061_out0;
wire  [3:0] v$_7116_out1;
wire  [3:0] v$_7117_out1;
wire  [3:0] v$_8687_out0;
wire  [3:0] v$_8688_out0;
wire  [3:0] v$_8689_out0;
wire  [3:0] v$_8690_out0;
wire  [4:0] v$0B00001_10554_out0;
wire  [4:0] v$0B00001_10555_out0;
wire  [4:0] v$A7_2719_out0;
wire  [4:0] v$A7_2720_out0;
wire  [4:0] v$B_3946_out0;
wire  [4:0] v$B_3947_out0;
wire  [4:0] v$C10_11248_out0;
wire  [4:0] v$C10_11249_out0;
wire  [4:0] v$C14_10795_out0;
wire  [4:0] v$C14_10796_out0;
wire  [4:0] v$C1_10313_out0;
wire  [4:0] v$C1_10314_out0;
wire  [4:0] v$C1_10315_out0;
wire  [4:0] v$C1_10316_out0;
wire  [4:0] v$C4_2593_out0;
wire  [4:0] v$C4_2594_out0;
wire  [4:0] v$C8_2758_out0;
wire  [4:0] v$C8_2759_out0;
wire  [4:0] v$EXP$ANS_10487_out0;
wire  [4:0] v$EXP$ANS_10488_out0;
wire  [4:0] v$EXP$ANS_10860_out0;
wire  [4:0] v$EXP$ANS_10861_out0;
wire  [4:0] v$EXP$ANS_11059_out0;
wire  [4:0] v$EXP$ANS_11060_out0;
wire  [4:0] v$EXP$ANS_13748_out0;
wire  [4:0] v$EXP$ANS_13749_out0;
wire  [4:0] v$EXP$ANS_2008_out0;
wire  [4:0] v$EXP$ANS_2009_out0;
wire  [4:0] v$EXP$PRE$ANS_10765_out0;
wire  [4:0] v$EXP$PRE$ANS_10766_out0;
wire  [4:0] v$EXP$RD_5855_out0;
wire  [4:0] v$EXP$RD_5856_out0;
wire  [4:0] v$EXP$RM_4743_out0;
wire  [4:0] v$EXP$RM_4744_out0;
wire  [4:0] v$EXP_2441_out0;
wire  [4:0] v$EXP_2442_out0;
wire  [4:0] v$EXP_2907_out0;
wire  [4:0] v$EXP_2908_out0;
wire  [4:0] v$K_2636_out0;
wire  [4:0] v$K_2637_out0;
wire  [4:0] v$K_5792_out0;
wire  [4:0] v$K_5793_out0;
wire  [4:0] v$MUX11_86_out0;
wire  [4:0] v$MUX11_87_out0;
wire  [4:0] v$MUX12_13783_out0;
wire  [4:0] v$MUX12_13784_out0;
wire  [4:0] v$MUX13_13647_out0;
wire  [4:0] v$MUX13_13648_out0;
wire  [4:0] v$MUX4_275_out0;
wire  [4:0] v$MUX4_276_out0;
wire  [4:0] v$MUX7_4481_out0;
wire  [4:0] v$MUX7_4482_out0;
wire  [4:0] v$OP2$EXP_10383_out0;
wire  [4:0] v$OP2$EXP_10384_out0;
wire  [4:0] v$OP2$EXP_2548_out0;
wire  [4:0] v$OP2$EXP_2549_out0;
wire  [4:0] v$OP2$EXP_536_out0;
wire  [4:0] v$OP2$EXP_537_out0;
wire  [4:0] v$RD$EXP_2601_out0;
wire  [4:0] v$RD$EXP_2602_out0;
wire  [4:0] v$RD$EXP_3951_out0;
wire  [4:0] v$RD$EXP_3952_out0;
wire  [4:0] v$RD$EXP_8846_out0;
wire  [4:0] v$RD$EXP_8847_out0;
wire  [4:0] v$SEL1_2917_out0;
wire  [4:0] v$SEL1_2918_out0;
wire  [4:0] v$SEL2_13327_out0;
wire  [4:0] v$SEL2_13328_out0;
wire  [4:0] v$SEL3_390_out0;
wire  [4:0] v$SEL3_391_out0;
wire  [4:0] v$SEL4_5790_out0;
wire  [4:0] v$SEL4_5791_out0;
wire  [4:0] v$SHIFT$AMOUNT_226_out0;
wire  [4:0] v$SHIFT$AMOUNT_227_out0;
wire  [4:0] v$SHIFT$AMOUNT_4715_out0;
wire  [4:0] v$SHIFT$AMOUNT_4716_out0;
wire  [4:0] v$_13518_out0;
wire  [4:0] v$_13519_out0;
wire  [4:0] v$_13520_out0;
wire  [4:0] v$_13521_out0;
wire  [4:0] v$_13522_out0;
wire  [4:0] v$_13523_out0;
wire  [4:0] v$_13524_out0;
wire  [4:0] v$_13525_out0;
wire  [4:0] v$_13526_out0;
wire  [4:0] v$_13527_out0;
wire  [4:0] v$_13528_out0;
wire  [4:0] v$_13529_out0;
wire  [4:0] v$_13530_out0;
wire  [4:0] v$_13531_out0;
wire  [4:0] v$_13532_out0;
wire  [4:0] v$_13533_out0;
wire  [4:0] v$_13534_out0;
wire  [4:0] v$_13535_out0;
wire  [4:0] v$_13536_out0;
wire  [4:0] v$_13537_out0;
wire  [4:0] v$_13538_out0;
wire  [4:0] v$_13539_out0;
wire  [4:0] v$_13540_out0;
wire  [4:0] v$_13541_out0;
wire  [4:0] v$_13542_out0;
wire  [4:0] v$_13543_out0;
wire  [4:0] v$_13544_out0;
wire  [4:0] v$_13545_out0;
wire  [4:0] v$_13546_out0;
wire  [4:0] v$_13547_out0;
wire  [4:0] v$_2392_out0;
wire  [4:0] v$_2393_out0;
wire  [4:0] v$_2846_out0;
wire  [4:0] v$_2847_out0;
wire  [4:0] v$_3251_out0;
wire  [4:0] v$_3252_out0;
wire  [4:0] v$_3253_out0;
wire  [4:0] v$_3254_out0;
wire  [4:0] v$_5849_out0;
wire  [4:0] v$_5850_out0;
wire  [5:0] v$A4_13603_out0;
wire  [5:0] v$A4_13604_out0;
wire  [5:0] v$A5_2638_out0;
wire  [5:0] v$A5_2639_out0;
wire  [5:0] v$A6_3957_out0;
wire  [5:0] v$A6_3958_out0;
wire  [5:0] v$C11_13765_out0;
wire  [5:0] v$C11_13766_out0;
wire  [5:0] v$C12_2113_out0;
wire  [5:0] v$C12_2114_out0;
wire  [5:0] v$C13_405_out0;
wire  [5:0] v$C13_406_out0;
wire  [5:0] v$C9_11159_out0;
wire  [5:0] v$C9_11160_out0;
wire  [5:0] v$EXP$SUM_5844_out0;
wire  [5:0] v$EXP$SUM_5845_out0;
wire  [5:0] v$MUX10_10395_out0;
wire  [5:0] v$MUX10_10396_out0;
wire  [5:0] v$MUX8_4587_out0;
wire  [5:0] v$MUX8_4588_out0;
wire  [5:0] v$MUX9_13486_out0;
wire  [5:0] v$MUX9_13487_out0;
wire  [5:0] v$NEG1_6921_out0;
wire  [5:0] v$NEG1_6922_out0;
wire  [5:0] v$NOTUSED_2698_out0;
wire  [5:0] v$NOTUSED_2699_out0;
wire  [5:0] v$XOR3_2546_out0;
wire  [5:0] v$XOR3_2547_out0;
wire  [5:0] v$XOR4_6960_out0;
wire  [5:0] v$XOR4_6961_out0;
wire  [5:0] v$_10262_out0;
wire  [5:0] v$_10263_out0;
wire  [5:0] v$_10298_out0;
wire  [5:0] v$_10299_out0;
wire  [5:0] v$_10300_out0;
wire  [5:0] v$_10301_out0;
wire  [5:0] v$_10490_out0;
wire  [5:0] v$_10491_out0;
wire  [5:0] v$_10858_out0;
wire  [5:0] v$_10859_out0;
wire  [5:0] v$_2610_out0;
wire  [5:0] v$_2611_out0;
wire  [5:0] v$_3311_out0;
wire  [5:0] v$_3312_out0;
wire  [5:0] v$_3313_out0;
wire  [5:0] v$_3314_out0;
wire  [5:0] v$_3315_out0;
wire  [5:0] v$_3316_out0;
wire  [5:0] v$_3317_out0;
wire  [5:0] v$_3318_out0;
wire  [5:0] v$_3319_out0;
wire  [5:0] v$_3320_out0;
wire  [5:0] v$_3321_out0;
wire  [5:0] v$_3322_out0;
wire  [5:0] v$_3323_out0;
wire  [5:0] v$_3324_out0;
wire  [5:0] v$_3325_out0;
wire  [5:0] v$_3326_out0;
wire  [5:0] v$_3327_out0;
wire  [5:0] v$_3328_out0;
wire  [5:0] v$_3329_out0;
wire  [5:0] v$_3330_out0;
wire  [5:0] v$_3331_out0;
wire  [5:0] v$_3332_out0;
wire  [5:0] v$_3333_out0;
wire  [5:0] v$_3334_out0;
wire  [5:0] v$_3335_out0;
wire  [5:0] v$_3336_out0;
wire  [5:0] v$_3337_out0;
wire  [5:0] v$_3338_out0;
wire  [5:0] v$_3339_out0;
wire  [5:0] v$_3340_out0;
wire  [5:0] v$_3897_out1;
wire  [5:0] v$_3898_out1;
wire  [5:0] v$_56_out0;
wire  [5:0] v$_57_out0;
wire  [5:0] v$_96_out0;
wire  [5:0] v$_97_out0;
wire  [6:0] v$_119_out0;
wire  [6:0] v$_120_out0;
wire  [6:0] v$_121_out0;
wire  [6:0] v$_122_out0;
wire  [6:0] v$_2959_out1;
wire  [6:0] v$_4703_out1;
wire  [6:0] v$_4704_out1;
wire  [6:0] v$_681_out0;
wire  [6:0] v$_682_out0;
wire  [6:0] v$_7062_out0;
wire  [6:0] v$_7063_out0;
wire  [6:0] v$_7147_out0;
wire  [6:0] v$_7148_out0;
wire  [6:0] v$_7149_out0;
wire  [6:0] v$_7150_out0;
wire  [6:0] v$_7151_out0;
wire  [6:0] v$_7152_out0;
wire  [6:0] v$_7153_out0;
wire  [6:0] v$_7154_out0;
wire  [6:0] v$_7155_out0;
wire  [6:0] v$_7156_out0;
wire  [6:0] v$_7157_out0;
wire  [6:0] v$_7158_out0;
wire  [6:0] v$_7159_out0;
wire  [6:0] v$_7160_out0;
wire  [6:0] v$_7161_out0;
wire  [6:0] v$_7162_out0;
wire  [6:0] v$_7163_out0;
wire  [6:0] v$_7164_out0;
wire  [6:0] v$_7165_out0;
wire  [6:0] v$_7166_out0;
wire  [6:0] v$_7167_out0;
wire  [6:0] v$_7168_out0;
wire  [6:0] v$_7169_out0;
wire  [6:0] v$_7170_out0;
wire  [6:0] v$_7171_out0;
wire  [6:0] v$_7172_out0;
wire  [6:0] v$_7173_out0;
wire  [6:0] v$_7174_out0;
wire  [6:0] v$_7175_out0;
wire  [6:0] v$_7176_out0;
wire  [6:0] v$_72_out0;
wire  [6:0] v$_73_out0;
wire  [7:0] v$BYTE$RECEIVED_13441_out0;
wire  [7:0] v$BYTE$RECEIVED_13796_out0;
wire  [7:0] v$BYTE$RECEIVED_2231_out0;
wire  [7:0] v$BYTE$RECEIVED_7101_out0;
wire  [7:0] v$BYTE$RECEIVED_7102_out0;
wire  [7:0] v$BYTE$RECEIVED_8819_out0;
wire  [7:0] v$BYTE$RECEIVED_8820_out0;
wire  [7:0] v$C1_10266_out0;
wire  [7:0] v$C1_10267_out0;
wire  [7:0] v$C1_13277_out0;
wire  [7:0] v$C1_13278_out0;
wire  [7:0] v$C1_13446_out0;
wire  [7:0] v$C1_13447_out0;
wire  [7:0] v$MUX1_13260_out0;
wire  [7:0] v$NOTUSED2_41_out0;
wire  [7:0] v$NOTUSED2_42_out0;
wire  [7:0] v$NOTUSED_10564_out0;
wire  [7:0] v$NOTUSED_10565_out0;
wire  [7:0] v$NOTUSED_683_out0;
wire  [7:0] v$NOTUSED_684_out0;
wire  [7:0] v$NOTUSED_68_out0;
wire  [7:0] v$NOTUSED_69_out0;
wire  [7:0] v$OUT_3037_out0;
wire  [7:0] v$RECEIVER$STREAM_564_out0;
wire  [7:0] v$RECEIVERSTREAM_7635_out0;
wire  [7:0] v$REGISTER$TRANSMIT$DATA_12241_out0;
wire  [7:0] v$TRANSIMISSION$DATA_10818_out0;
wire  [7:0] v$TRANSMISSION$DATA2_7014_out0;
wire  [7:0] v$TRANSMIT$DATA_76_out0;
wire  [7:0] v$_10376_out0;
wire  [7:0] v$_10868_out0;
wire  [7:0] v$_10869_out0;
wire  [7:0] v$_11132_out0;
wire  [7:0] v$_11132_out1;
wire  [7:0] v$_11133_out0;
wire  [7:0] v$_11133_out1;
wire  [7:0] v$_13790_out0;
wire  [7:0] v$_13791_out0;
wire  [7:0] v$_13792_out0;
wire  [7:0] v$_13793_out0;
wire  [7:0] v$_2425_out0;
wire  [7:0] v$_2437_out1;
wire  [7:0] v$_2438_out1;
wire  [7:0] v$_2582_out0;
wire  [7:0] v$_2582_out1;
wire  [7:0] v$_2583_out0;
wire  [7:0] v$_2583_out1;
wire  [7:0] v$_2680_out0;
wire  [7:0] v$_2681_out0;
wire  [7:0] v$_2684_out0;
wire  [7:0] v$_2685_out0;
wire  [7:0] v$_2686_out0;
wire  [7:0] v$_2687_out0;
wire  [7:0] v$_3040_out0;
wire  [7:0] v$_3125_out0;
wire  [7:0] v$_3125_out1;
wire  [7:0] v$_3126_out0;
wire  [7:0] v$_3126_out1;
wire  [7:0] v$_4449_out0;
wire  [7:0] v$_4450_out0;
wire  [7:0] v$_4451_out0;
wire  [7:0] v$_4452_out0;
wire  [7:0] v$_4749_out0;
wire  [7:0] v$_4750_out0;
wire  [7:0] v$_4751_out0;
wire  [7:0] v$_4752_out0;
wire  [7:0] v$_4753_out0;
wire  [7:0] v$_4754_out0;
wire  [7:0] v$_4755_out0;
wire  [7:0] v$_4756_out0;
wire  [7:0] v$_4757_out0;
wire  [7:0] v$_4758_out0;
wire  [7:0] v$_4759_out0;
wire  [7:0] v$_4760_out0;
wire  [7:0] v$_4761_out0;
wire  [7:0] v$_4762_out0;
wire  [7:0] v$_4763_out0;
wire  [7:0] v$_4764_out0;
wire  [7:0] v$_4765_out0;
wire  [7:0] v$_4766_out0;
wire  [7:0] v$_4767_out0;
wire  [7:0] v$_4768_out0;
wire  [7:0] v$_4769_out0;
wire  [7:0] v$_4770_out0;
wire  [7:0] v$_4771_out0;
wire  [7:0] v$_4772_out0;
wire  [7:0] v$_4773_out0;
wire  [7:0] v$_4774_out0;
wire  [7:0] v$_4775_out0;
wire  [7:0] v$_4776_out0;
wire  [7:0] v$_4777_out0;
wire  [7:0] v$_4778_out0;
wire  [7:0] v$_636_out0;
wire  [7:0] v$_637_out0;
wire  [7:0] v$_8673_out0;
wire  [7:0] v$_8673_out1;
wire  [7:0] v$_8674_out0;
wire  [7:0] v$_8674_out1;
wire  [7:0] v$_8681_out0;
wire  [7:0] v$_8682_out0;
wire  [7:0] v$split_3196_out0;
wire  [7:0] v$split_3196_out1;
wire  [8:0] v$SEL6_3991_out0;
wire  [8:0] v$SEL6_3992_out0;
wire  [8:0] v$_13550_out1;
wire  [8:0] v$_13551_out1;
wire  [8:0] v$_2838_out0;
wire  [8:0] v$_2839_out0;
wire  [8:0] v$_43_out0;
wire  [8:0] v$_44_out0;
wire  [8:0] v$_4526_out0;
wire  [8:0] v$_4527_out0;
wire  [8:0] v$_464_out0;
wire  [8:0] v$_465_out0;
wire  [8:0] v$_466_out0;
wire  [8:0] v$_467_out0;
wire  [8:0] v$_6926_out0;
wire  [8:0] v$_6927_out0;
wire  [8:0] v$_6928_out0;
wire  [8:0] v$_6929_out0;
wire  [8:0] v$_6930_out0;
wire  [8:0] v$_6931_out0;
wire  [8:0] v$_6932_out0;
wire  [8:0] v$_6933_out0;
wire  [8:0] v$_6934_out0;
wire  [8:0] v$_6935_out0;
wire  [8:0] v$_6936_out0;
wire  [8:0] v$_6937_out0;
wire  [8:0] v$_6938_out0;
wire  [8:0] v$_6939_out0;
wire  [8:0] v$_6940_out0;
wire  [8:0] v$_6941_out0;
wire  [8:0] v$_6942_out0;
wire  [8:0] v$_6943_out0;
wire  [8:0] v$_6944_out0;
wire  [8:0] v$_6945_out0;
wire  [8:0] v$_6946_out0;
wire  [8:0] v$_6947_out0;
wire  [8:0] v$_6948_out0;
wire  [8:0] v$_6949_out0;
wire  [8:0] v$_6950_out0;
wire  [8:0] v$_6951_out0;
wire  [8:0] v$_6952_out0;
wire  [8:0] v$_6953_out0;
wire  [8:0] v$_6954_out0;
wire  [8:0] v$_6955_out0;
wire  [8:0] v$_7704_out0;
wire  [8:0] v$_7705_out0;
wire  [9:0] v$MUX4_10357_out0;
wire  [9:0] v$MUX4_10358_out0;
wire  [9:0] v$MUX6_10350_out0;
wire  [9:0] v$MUX6_10351_out0;
wire  [9:0] v$OP2$SIG_13301_out0;
wire  [9:0] v$OP2$SIG_13302_out0;
wire  [9:0] v$RD$SIG_1769_out0;
wire  [9:0] v$RD$SIG_1770_out0;
wire  [9:0] v$SEL4_11225_out0;
wire  [9:0] v$SEL4_11226_out0;
wire  [9:0] v$SEL5_8767_out0;
wire  [9:0] v$SEL5_8768_out0;
wire  [9:0] v$SEL6_103_out0;
wire  [9:0] v$SEL6_104_out0;
wire  [9:0] v$SEL9_13753_out0;
wire  [9:0] v$SEL9_13754_out0;
wire  [9:0] v$SIG$ANS_10296_out0;
wire  [9:0] v$SIG$ANS_10297_out0;
wire  [9:0] v$SIG$ANS_2335_out0;
wire  [9:0] v$SIG$ANS_2336_out0;
wire  [9:0] v$SIG$ANS_3276_out0;
wire  [9:0] v$SIG$ANS_3277_out0;
wire  [9:0] v$SIG$ANS_439_out0;
wire  [9:0] v$SIG$ANS_440_out0;
wire  [9:0] v$SIG$RD_11298_out0;
wire  [9:0] v$SIG$RD_11299_out0;
wire  [9:0] v$SIG$RM_1767_out0;
wire  [9:0] v$SIG$RM_1768_out0;
wire  [9:0] v$_10775_out0;
wire  [9:0] v$_10776_out0;
wire  [9:0] v$_10806_out0;
wire  [9:0] v$_10807_out0;
wire  [9:0] v$_2649_out0;
wire  [9:0] v$_2650_out0;
wire  [9:0] v$_3897_out0;
wire  [9:0] v$_3898_out0;
wire  [9:0] v$_3907_out1;
wire  [9:0] v$_3908_out1;
wire  [9:0] v$_422_out0;
wire  [9:0] v$_423_out0;
wire  [9:0] v$_424_out0;
wire  [9:0] v$_425_out0;
wire  [9:0] v$_5802_out0;
wire  [9:0] v$_5803_out0;
wire  [9:0] v$_5804_out0;
wire  [9:0] v$_5805_out0;
wire  [9:0] v$_5806_out0;
wire  [9:0] v$_5807_out0;
wire  [9:0] v$_5808_out0;
wire  [9:0] v$_5809_out0;
wire  [9:0] v$_5810_out0;
wire  [9:0] v$_5811_out0;
wire  [9:0] v$_5812_out0;
wire  [9:0] v$_5813_out0;
wire  [9:0] v$_5814_out0;
wire  [9:0] v$_5815_out0;
wire  [9:0] v$_5816_out0;
wire  [9:0] v$_5817_out0;
wire  [9:0] v$_5818_out0;
wire  [9:0] v$_5819_out0;
wire  [9:0] v$_5820_out0;
wire  [9:0] v$_5821_out0;
wire  [9:0] v$_5822_out0;
wire  [9:0] v$_5823_out0;
wire  [9:0] v$_5824_out0;
wire  [9:0] v$_5825_out0;
wire  [9:0] v$_5826_out0;
wire  [9:0] v$_5827_out0;
wire  [9:0] v$_5828_out0;
wire  [9:0] v$_5829_out0;
wire  [9:0] v$_5830_out0;
wire  [9:0] v$_5831_out0;
wire  [9:0] v$_8677_out0;
wire  [9:0] v$_8678_out0;
wire v$0_10706_out0;
wire v$0_10707_out0;
wire v$0_3022_out0;
wire v$0_3023_out0;
wire v$1_3817_out0;
wire v$1_3818_out0;
wire v$2_1763_out0;
wire v$2_1764_out0;
wire v$2_7072_out0;
wire v$3_13619_out0;
wire v$3_13620_out0;
wire v$9_13623_out0;
wire v$9_13624_out0;
wire v$9_13625_out0;
wire v$9_13626_out0;
wire v$9_1700_out0;
wire v$9_1701_out0;
wire v$9_1702_out0;
wire v$9_1703_out0;
wire v$9_417_out0;
wire v$A1_11043_out1;
wire v$A1_3174_out1;
wire v$A1_3175_out1;
wire v$A1_3855_out1;
wire v$A1_3856_out1;
wire v$A1_7019_out1;
wire v$A1_7020_out1;
wire v$A4_11227_out1;
wire v$A4_11228_out1;
wire v$A4_13603_out1;
wire v$A4_13604_out1;
wire v$A5_1901_out1;
wire v$A5_1902_out1;
wire v$A5_2638_out1;
wire v$A5_2639_out1;
wire v$A6_10463_out1;
wire v$A6_10464_out1;
wire v$A6_3957_out1;
wire v$A6_3958_out1;
wire v$A7_2719_out1;
wire v$A7_2720_out1;
wire v$A8_11155_out1;
wire v$A8_11156_out1;
wire v$ADC_10393_out0;
wire v$ADC_10394_out0;
wire v$ADC_13614_out0;
wire v$ADC_13615_out0;
wire v$ADC_1821_out0;
wire v$ADC_1822_out0;
wire v$ADD_11193_out0;
wire v$ADD_11194_out0;
wire v$ADD_4455_out0;
wire v$ADD_4456_out0;
wire v$AND_13556_out0;
wire v$AND_13557_out0;
wire v$AND_3858_out0;
wire v$AND_3859_out0;
wire v$ASR_10366_out0;
wire v$ASR_10367_out0;
wire v$ASR_10566_out0;
wire v$ASR_10567_out0;
wire v$ASR_13713_out0;
wire v$ASR_13714_out0;
wire v$ASR_8754_out0;
wire v$ASR_8755_out0;
wire v$BIT$IN1_3209_out0;
wire v$BIT$OUT_10705_out0;
wire v$BIT$OUT_13326_out0;
wire v$BIT$OUT_2015_out0;
wire v$BIT$STREAM$IN_13_out0;
wire v$BIT10_7009_out0;
wire v$BIT10_7010_out0;
wire v$BIT_2328_out0;
wire v$BIT_383_out0;
wire v$BIT_6918_out0;
wire v$BYTE$COMP$10_13611_out0;
wire v$BYTE$COMP$11_1163_out0;
wire v$BYTE$COMP$1_8743_out0;
wire v$BYTE$COMP1_3262_out0;
wire v$BYTE$COMP1_3263_out0;
wire v$BYTE$COMP1_9796_out0;
wire v$BYTE$COMP1_9797_out0;
wire v$BYTE$READY_10558_out0;
wire v$BYTE$READY_10559_out0;
wire v$BYTE$READY_11172_out0;
wire v$BYTE$READY_11173_out0;
wire v$BYTE$READY_13255_out0;
wire v$BYTE$READY_2852_out0;
wire v$BYTE$READY_2853_out0;
wire v$BYTE$READY_7021_out0;
wire v$BYTE$READY_7022_out0;
wire v$BYTE1$comp1_2443_out0;
wire v$BYTE1$comp1_2444_out0;
wire v$BYTE2$COMP8_7695_out0;
wire v$BYTE2$COMP8_7696_out0;
wire v$BYTERECEIVED_11197_out0;
wire v$C10_1819_out0;
wire v$C10_1820_out0;
wire v$C12_1151_out0;
wire v$C12_1152_out0;
wire v$C14_1674_out0;
wire v$C14_1675_out0;
wire v$C1_10259_out0;
wire v$C1_10789_out0;
wire v$C1_10790_out0;
wire v$C1_436_out0;
wire v$C1_604_out0;
wire v$C1_605_out0;
wire v$C1_8815_out0;
wire v$C1_8816_out0;
wire v$C3_2764_out0;
wire v$C3_4741_out0;
wire v$C3_4742_out0;
wire v$C4_10619_out0;
wire v$C4_90_out0;
wire v$C5_11031_out0;
wire v$C5_13267_out0;
wire v$C6_10317_out0;
wire v$C6_10318_out0;
wire v$C6_1732_out0;
wire v$C7_2271_out0;
wire v$C7_2272_out0;
wire v$C7_3222_out0;
wire v$C9_3029_out0;
wire v$C9_3030_out0;
wire v$CARRY_4862_out0;
wire v$CARRY_4863_out0;
wire v$CARRY_4864_out0;
wire v$CARRY_4865_out0;
wire v$CARRY_4866_out0;
wire v$CARRY_4867_out0;
wire v$CARRY_4868_out0;
wire v$CARRY_4869_out0;
wire v$CARRY_4870_out0;
wire v$CARRY_4871_out0;
wire v$CARRY_4872_out0;
wire v$CARRY_4873_out0;
wire v$CARRY_4874_out0;
wire v$CARRY_4875_out0;
wire v$CARRY_4876_out0;
wire v$CARRY_4877_out0;
wire v$CARRY_4878_out0;
wire v$CARRY_4879_out0;
wire v$CARRY_4880_out0;
wire v$CARRY_4881_out0;
wire v$CARRY_4882_out0;
wire v$CARRY_4883_out0;
wire v$CARRY_4884_out0;
wire v$CARRY_4885_out0;
wire v$CARRY_4886_out0;
wire v$CARRY_4887_out0;
wire v$CARRY_4888_out0;
wire v$CARRY_4889_out0;
wire v$CARRY_4890_out0;
wire v$CARRY_4891_out0;
wire v$CARRY_4892_out0;
wire v$CARRY_4893_out0;
wire v$CARRY_4894_out0;
wire v$CARRY_4895_out0;
wire v$CARRY_4896_out0;
wire v$CARRY_4897_out0;
wire v$CARRY_4898_out0;
wire v$CARRY_4899_out0;
wire v$CARRY_4900_out0;
wire v$CARRY_4901_out0;
wire v$CARRY_4902_out0;
wire v$CARRY_4903_out0;
wire v$CARRY_4904_out0;
wire v$CARRY_4905_out0;
wire v$CARRY_4906_out0;
wire v$CARRY_4907_out0;
wire v$CARRY_4908_out0;
wire v$CARRY_4909_out0;
wire v$CARRY_4910_out0;
wire v$CARRY_4911_out0;
wire v$CARRY_4912_out0;
wire v$CARRY_4913_out0;
wire v$CARRY_4914_out0;
wire v$CARRY_4915_out0;
wire v$CARRY_4916_out0;
wire v$CARRY_4917_out0;
wire v$CARRY_4918_out0;
wire v$CARRY_4919_out0;
wire v$CARRY_4920_out0;
wire v$CARRY_4921_out0;
wire v$CARRY_4922_out0;
wire v$CARRY_4923_out0;
wire v$CARRY_4924_out0;
wire v$CARRY_4925_out0;
wire v$CARRY_4926_out0;
wire v$CARRY_4927_out0;
wire v$CARRY_4928_out0;
wire v$CARRY_4929_out0;
wire v$CARRY_4930_out0;
wire v$CARRY_4931_out0;
wire v$CARRY_4932_out0;
wire v$CARRY_4933_out0;
wire v$CARRY_4934_out0;
wire v$CARRY_4935_out0;
wire v$CARRY_4936_out0;
wire v$CARRY_4937_out0;
wire v$CARRY_4938_out0;
wire v$CARRY_4939_out0;
wire v$CARRY_4940_out0;
wire v$CARRY_4941_out0;
wire v$CARRY_4942_out0;
wire v$CARRY_4943_out0;
wire v$CARRY_4944_out0;
wire v$CARRY_4945_out0;
wire v$CARRY_4946_out0;
wire v$CARRY_4947_out0;
wire v$CARRY_4948_out0;
wire v$CARRY_4949_out0;
wire v$CARRY_4950_out0;
wire v$CARRY_4951_out0;
wire v$CARRY_4952_out0;
wire v$CARRY_4953_out0;
wire v$CARRY_4954_out0;
wire v$CARRY_4955_out0;
wire v$CARRY_4956_out0;
wire v$CARRY_4957_out0;
wire v$CARRY_4958_out0;
wire v$CARRY_4959_out0;
wire v$CARRY_4960_out0;
wire v$CARRY_4961_out0;
wire v$CARRY_4962_out0;
wire v$CARRY_4963_out0;
wire v$CARRY_4964_out0;
wire v$CARRY_4965_out0;
wire v$CARRY_4966_out0;
wire v$CARRY_4967_out0;
wire v$CARRY_4968_out0;
wire v$CARRY_4969_out0;
wire v$CARRY_4970_out0;
wire v$CARRY_4971_out0;
wire v$CARRY_4972_out0;
wire v$CARRY_4973_out0;
wire v$CARRY_4974_out0;
wire v$CARRY_4975_out0;
wire v$CARRY_4976_out0;
wire v$CARRY_4977_out0;
wire v$CARRY_4978_out0;
wire v$CARRY_4979_out0;
wire v$CARRY_4980_out0;
wire v$CARRY_4981_out0;
wire v$CARRY_4982_out0;
wire v$CARRY_4983_out0;
wire v$CARRY_4984_out0;
wire v$CARRY_4985_out0;
wire v$CARRY_4986_out0;
wire v$CARRY_4987_out0;
wire v$CARRY_4988_out0;
wire v$CARRY_4989_out0;
wire v$CARRY_4990_out0;
wire v$CARRY_4991_out0;
wire v$CARRY_4992_out0;
wire v$CARRY_4993_out0;
wire v$CARRY_4994_out0;
wire v$CARRY_4995_out0;
wire v$CARRY_4996_out0;
wire v$CARRY_4997_out0;
wire v$CARRY_4998_out0;
wire v$CARRY_4999_out0;
wire v$CARRY_5000_out0;
wire v$CARRY_5001_out0;
wire v$CARRY_5002_out0;
wire v$CARRY_5003_out0;
wire v$CARRY_5004_out0;
wire v$CARRY_5005_out0;
wire v$CARRY_5006_out0;
wire v$CARRY_5007_out0;
wire v$CARRY_5008_out0;
wire v$CARRY_5009_out0;
wire v$CARRY_5010_out0;
wire v$CARRY_5011_out0;
wire v$CARRY_5012_out0;
wire v$CARRY_5013_out0;
wire v$CARRY_5014_out0;
wire v$CARRY_5015_out0;
wire v$CARRY_5016_out0;
wire v$CARRY_5017_out0;
wire v$CARRY_5018_out0;
wire v$CARRY_5019_out0;
wire v$CARRY_5020_out0;
wire v$CARRY_5021_out0;
wire v$CARRY_5022_out0;
wire v$CARRY_5023_out0;
wire v$CARRY_5024_out0;
wire v$CARRY_5025_out0;
wire v$CARRY_5026_out0;
wire v$CARRY_5027_out0;
wire v$CARRY_5028_out0;
wire v$CARRY_5029_out0;
wire v$CARRY_5030_out0;
wire v$CARRY_5031_out0;
wire v$CARRY_5032_out0;
wire v$CARRY_5033_out0;
wire v$CARRY_5034_out0;
wire v$CARRY_5035_out0;
wire v$CARRY_5036_out0;
wire v$CARRY_5037_out0;
wire v$CARRY_5038_out0;
wire v$CARRY_5039_out0;
wire v$CARRY_5040_out0;
wire v$CARRY_5041_out0;
wire v$CARRY_5042_out0;
wire v$CARRY_5043_out0;
wire v$CARRY_5044_out0;
wire v$CARRY_5045_out0;
wire v$CARRY_5046_out0;
wire v$CARRY_5047_out0;
wire v$CARRY_5048_out0;
wire v$CARRY_5049_out0;
wire v$CARRY_5050_out0;
wire v$CARRY_5051_out0;
wire v$CARRY_5052_out0;
wire v$CARRY_5053_out0;
wire v$CARRY_5054_out0;
wire v$CARRY_5055_out0;
wire v$CARRY_5056_out0;
wire v$CARRY_5057_out0;
wire v$CARRY_5058_out0;
wire v$CARRY_5059_out0;
wire v$CARRY_5060_out0;
wire v$CARRY_5061_out0;
wire v$CARRY_5062_out0;
wire v$CARRY_5063_out0;
wire v$CARRY_5064_out0;
wire v$CARRY_5065_out0;
wire v$CARRY_5066_out0;
wire v$CARRY_5067_out0;
wire v$CARRY_5068_out0;
wire v$CARRY_5069_out0;
wire v$CARRY_5070_out0;
wire v$CARRY_5071_out0;
wire v$CARRY_5072_out0;
wire v$CARRY_5073_out0;
wire v$CARRY_5074_out0;
wire v$CARRY_5075_out0;
wire v$CARRY_5076_out0;
wire v$CARRY_5077_out0;
wire v$CARRY_5078_out0;
wire v$CARRY_5079_out0;
wire v$CARRY_5080_out0;
wire v$CARRY_5081_out0;
wire v$CARRY_5082_out0;
wire v$CARRY_5083_out0;
wire v$CARRY_5084_out0;
wire v$CARRY_5085_out0;
wire v$CARRY_5086_out0;
wire v$CARRY_5087_out0;
wire v$CARRY_5088_out0;
wire v$CARRY_5089_out0;
wire v$CARRY_5090_out0;
wire v$CARRY_5091_out0;
wire v$CARRY_5092_out0;
wire v$CARRY_5093_out0;
wire v$CARRY_5094_out0;
wire v$CARRY_5095_out0;
wire v$CARRY_5096_out0;
wire v$CARRY_5097_out0;
wire v$CARRY_5098_out0;
wire v$CARRY_5099_out0;
wire v$CARRY_5100_out0;
wire v$CARRY_5101_out0;
wire v$CARRY_5102_out0;
wire v$CARRY_5103_out0;
wire v$CARRY_5104_out0;
wire v$CARRY_5105_out0;
wire v$CARRY_5106_out0;
wire v$CARRY_5107_out0;
wire v$CARRY_5108_out0;
wire v$CARRY_5109_out0;
wire v$CARRY_5110_out0;
wire v$CARRY_5111_out0;
wire v$CARRY_5112_out0;
wire v$CARRY_5113_out0;
wire v$CARRY_5114_out0;
wire v$CARRY_5115_out0;
wire v$CARRY_5116_out0;
wire v$CARRY_5117_out0;
wire v$CARRY_5118_out0;
wire v$CARRY_5119_out0;
wire v$CARRY_5120_out0;
wire v$CARRY_5121_out0;
wire v$CARRY_5122_out0;
wire v$CARRY_5123_out0;
wire v$CARRY_5124_out0;
wire v$CARRY_5125_out0;
wire v$CARRY_5126_out0;
wire v$CARRY_5127_out0;
wire v$CARRY_5128_out0;
wire v$CARRY_5129_out0;
wire v$CARRY_5130_out0;
wire v$CARRY_5131_out0;
wire v$CARRY_5132_out0;
wire v$CARRY_5133_out0;
wire v$CARRY_5134_out0;
wire v$CARRY_5135_out0;
wire v$CARRY_5136_out0;
wire v$CARRY_5137_out0;
wire v$CARRY_5138_out0;
wire v$CARRY_5139_out0;
wire v$CARRY_5140_out0;
wire v$CARRY_5141_out0;
wire v$CARRY_5142_out0;
wire v$CARRY_5143_out0;
wire v$CARRY_5144_out0;
wire v$CARRY_5145_out0;
wire v$CARRY_5146_out0;
wire v$CARRY_5147_out0;
wire v$CARRY_5148_out0;
wire v$CARRY_5149_out0;
wire v$CARRY_5150_out0;
wire v$CARRY_5151_out0;
wire v$CARRY_5152_out0;
wire v$CARRY_5153_out0;
wire v$CARRY_5154_out0;
wire v$CARRY_5155_out0;
wire v$CARRY_5156_out0;
wire v$CARRY_5157_out0;
wire v$CARRY_5158_out0;
wire v$CARRY_5159_out0;
wire v$CARRY_5160_out0;
wire v$CARRY_5161_out0;
wire v$CARRY_5162_out0;
wire v$CARRY_5163_out0;
wire v$CARRY_5164_out0;
wire v$CARRY_5165_out0;
wire v$CARRY_5166_out0;
wire v$CARRY_5167_out0;
wire v$CARRY_5168_out0;
wire v$CARRY_5169_out0;
wire v$CARRY_5170_out0;
wire v$CARRY_5171_out0;
wire v$CARRY_5172_out0;
wire v$CARRY_5173_out0;
wire v$CARRY_5174_out0;
wire v$CARRY_5175_out0;
wire v$CARRY_5176_out0;
wire v$CARRY_5177_out0;
wire v$CARRY_5178_out0;
wire v$CARRY_5179_out0;
wire v$CARRY_5180_out0;
wire v$CARRY_5181_out0;
wire v$CARRY_5182_out0;
wire v$CARRY_5183_out0;
wire v$CARRY_5184_out0;
wire v$CARRY_5185_out0;
wire v$CARRY_5186_out0;
wire v$CARRY_5187_out0;
wire v$CARRY_5188_out0;
wire v$CARRY_5189_out0;
wire v$CARRY_5190_out0;
wire v$CARRY_5191_out0;
wire v$CARRY_5192_out0;
wire v$CARRY_5193_out0;
wire v$CARRY_5194_out0;
wire v$CARRY_5195_out0;
wire v$CARRY_5196_out0;
wire v$CARRY_5197_out0;
wire v$CARRY_5198_out0;
wire v$CARRY_5199_out0;
wire v$CARRY_5200_out0;
wire v$CARRY_5201_out0;
wire v$CARRY_5202_out0;
wire v$CARRY_5203_out0;
wire v$CARRY_5204_out0;
wire v$CARRY_5205_out0;
wire v$CARRY_5206_out0;
wire v$CARRY_5207_out0;
wire v$CARRY_5208_out0;
wire v$CARRY_5209_out0;
wire v$CARRY_5210_out0;
wire v$CARRY_5211_out0;
wire v$CARRY_5212_out0;
wire v$CARRY_5213_out0;
wire v$CARRY_5214_out0;
wire v$CARRY_5215_out0;
wire v$CARRY_5216_out0;
wire v$CARRY_5217_out0;
wire v$CARRY_5218_out0;
wire v$CARRY_5219_out0;
wire v$CARRY_5220_out0;
wire v$CARRY_5221_out0;
wire v$CARRY_5222_out0;
wire v$CARRY_5223_out0;
wire v$CARRY_5224_out0;
wire v$CARRY_5225_out0;
wire v$CARRY_5226_out0;
wire v$CARRY_5227_out0;
wire v$CARRY_5228_out0;
wire v$CARRY_5229_out0;
wire v$CARRY_5230_out0;
wire v$CARRY_5231_out0;
wire v$CARRY_5232_out0;
wire v$CARRY_5233_out0;
wire v$CARRY_5234_out0;
wire v$CARRY_5235_out0;
wire v$CARRY_5236_out0;
wire v$CARRY_5237_out0;
wire v$CARRY_5238_out0;
wire v$CARRY_5239_out0;
wire v$CARRY_5240_out0;
wire v$CARRY_5241_out0;
wire v$CARRY_5242_out0;
wire v$CARRY_5243_out0;
wire v$CARRY_5244_out0;
wire v$CARRY_5245_out0;
wire v$CARRY_5246_out0;
wire v$CARRY_5247_out0;
wire v$CARRY_5248_out0;
wire v$CARRY_5249_out0;
wire v$CARRY_5250_out0;
wire v$CARRY_5251_out0;
wire v$CARRY_5252_out0;
wire v$CARRY_5253_out0;
wire v$CARRY_5254_out0;
wire v$CARRY_5255_out0;
wire v$CARRY_5256_out0;
wire v$CARRY_5257_out0;
wire v$CARRY_5258_out0;
wire v$CARRY_5259_out0;
wire v$CARRY_5260_out0;
wire v$CARRY_5261_out0;
wire v$CARRY_5262_out0;
wire v$CARRY_5263_out0;
wire v$CARRY_5264_out0;
wire v$CARRY_5265_out0;
wire v$CARRY_5266_out0;
wire v$CARRY_5267_out0;
wire v$CARRY_5268_out0;
wire v$CARRY_5269_out0;
wire v$CARRY_5270_out0;
wire v$CARRY_5271_out0;
wire v$CARRY_5272_out0;
wire v$CARRY_5273_out0;
wire v$CARRY_5274_out0;
wire v$CARRY_5275_out0;
wire v$CARRY_5276_out0;
wire v$CARRY_5277_out0;
wire v$CARRY_5278_out0;
wire v$CARRY_5279_out0;
wire v$CARRY_5280_out0;
wire v$CARRY_5281_out0;
wire v$CARRY_5282_out0;
wire v$CARRY_5283_out0;
wire v$CARRY_5284_out0;
wire v$CARRY_5285_out0;
wire v$CARRY_5286_out0;
wire v$CARRY_5287_out0;
wire v$CARRY_5288_out0;
wire v$CARRY_5289_out0;
wire v$CARRY_5290_out0;
wire v$CARRY_5291_out0;
wire v$CARRY_5292_out0;
wire v$CARRY_5293_out0;
wire v$CARRY_5294_out0;
wire v$CARRY_5295_out0;
wire v$CARRY_5296_out0;
wire v$CARRY_5297_out0;
wire v$CARRY_5298_out0;
wire v$CARRY_5299_out0;
wire v$CARRY_5300_out0;
wire v$CARRY_5301_out0;
wire v$CARRY_5302_out0;
wire v$CARRY_5303_out0;
wire v$CARRY_5304_out0;
wire v$CARRY_5305_out0;
wire v$CARRY_5306_out0;
wire v$CARRY_5307_out0;
wire v$CARRY_5308_out0;
wire v$CARRY_5309_out0;
wire v$CARRY_5310_out0;
wire v$CARRY_5311_out0;
wire v$CARRY_5312_out0;
wire v$CARRY_5313_out0;
wire v$CARRY_5314_out0;
wire v$CARRY_5315_out0;
wire v$CARRY_5316_out0;
wire v$CARRY_5317_out0;
wire v$CARRY_5318_out0;
wire v$CARRY_5319_out0;
wire v$CARRY_5320_out0;
wire v$CARRY_5321_out0;
wire v$CARRY_5322_out0;
wire v$CARRY_5323_out0;
wire v$CARRY_5324_out0;
wire v$CARRY_5325_out0;
wire v$CARRY_5326_out0;
wire v$CARRY_5327_out0;
wire v$CARRY_5328_out0;
wire v$CARRY_5329_out0;
wire v$CARRY_5330_out0;
wire v$CARRY_5331_out0;
wire v$CARRY_5332_out0;
wire v$CARRY_5333_out0;
wire v$CARRY_5334_out0;
wire v$CARRY_5335_out0;
wire v$CARRY_5336_out0;
wire v$CARRY_5337_out0;
wire v$CARRY_5338_out0;
wire v$CARRY_5339_out0;
wire v$CARRY_5340_out0;
wire v$CARRY_5341_out0;
wire v$CARRY_5342_out0;
wire v$CARRY_5343_out0;
wire v$CARRY_5344_out0;
wire v$CARRY_5345_out0;
wire v$CARRY_5346_out0;
wire v$CARRY_5347_out0;
wire v$CARRY_5348_out0;
wire v$CARRY_5349_out0;
wire v$CARRY_5350_out0;
wire v$CARRY_5351_out0;
wire v$CARRY_5352_out0;
wire v$CARRY_5353_out0;
wire v$CARRY_5354_out0;
wire v$CARRY_5355_out0;
wire v$CARRY_5356_out0;
wire v$CARRY_5357_out0;
wire v$CARRY_5358_out0;
wire v$CARRY_5359_out0;
wire v$CARRY_5360_out0;
wire v$CARRY_5361_out0;
wire v$CARRY_5362_out0;
wire v$CARRY_5363_out0;
wire v$CARRY_5364_out0;
wire v$CARRY_5365_out0;
wire v$CARRY_5366_out0;
wire v$CARRY_5367_out0;
wire v$CARRY_5368_out0;
wire v$CARRY_5369_out0;
wire v$CARRY_5370_out0;
wire v$CARRY_5371_out0;
wire v$CARRY_5372_out0;
wire v$CARRY_5373_out0;
wire v$CARRY_5374_out0;
wire v$CARRY_5375_out0;
wire v$CARRY_5376_out0;
wire v$CARRY_5377_out0;
wire v$CARRY_5378_out0;
wire v$CARRY_5379_out0;
wire v$CARRY_5380_out0;
wire v$CARRY_5381_out0;
wire v$CARRY_5382_out0;
wire v$CARRY_5383_out0;
wire v$CARRY_5384_out0;
wire v$CARRY_5385_out0;
wire v$CARRY_5386_out0;
wire v$CARRY_5387_out0;
wire v$CARRY_5388_out0;
wire v$CARRY_5389_out0;
wire v$CARRY_5390_out0;
wire v$CARRY_5391_out0;
wire v$CARRY_5392_out0;
wire v$CARRY_5393_out0;
wire v$CARRY_5394_out0;
wire v$CARRY_5395_out0;
wire v$CARRY_5396_out0;
wire v$CARRY_5397_out0;
wire v$CARRY_5398_out0;
wire v$CARRY_5399_out0;
wire v$CARRY_5400_out0;
wire v$CARRY_5401_out0;
wire v$CARRY_5402_out0;
wire v$CARRY_5403_out0;
wire v$CARRY_5404_out0;
wire v$CARRY_5405_out0;
wire v$CARRY_5406_out0;
wire v$CARRY_5407_out0;
wire v$CARRY_5408_out0;
wire v$CARRY_5409_out0;
wire v$CARRY_5410_out0;
wire v$CARRY_5411_out0;
wire v$CARRY_5412_out0;
wire v$CARRY_5413_out0;
wire v$CARRY_5414_out0;
wire v$CARRY_5415_out0;
wire v$CARRY_5416_out0;
wire v$CARRY_5417_out0;
wire v$CARRY_5418_out0;
wire v$CARRY_5419_out0;
wire v$CARRY_5420_out0;
wire v$CARRY_5421_out0;
wire v$CARRY_5422_out0;
wire v$CARRY_5423_out0;
wire v$CARRY_5424_out0;
wire v$CARRY_5425_out0;
wire v$CARRY_5426_out0;
wire v$CARRY_5427_out0;
wire v$CARRY_5428_out0;
wire v$CARRY_5429_out0;
wire v$CARRY_5430_out0;
wire v$CARRY_5431_out0;
wire v$CARRY_5432_out0;
wire v$CARRY_5433_out0;
wire v$CARRY_5434_out0;
wire v$CARRY_5435_out0;
wire v$CARRY_5436_out0;
wire v$CARRY_5437_out0;
wire v$CARRY_5438_out0;
wire v$CARRY_5439_out0;
wire v$CARRY_5440_out0;
wire v$CARRY_5441_out0;
wire v$CARRY_5442_out0;
wire v$CARRY_5443_out0;
wire v$CARRY_5444_out0;
wire v$CARRY_5445_out0;
wire v$CARRY_5446_out0;
wire v$CARRY_5447_out0;
wire v$CARRY_5448_out0;
wire v$CARRY_5449_out0;
wire v$CARRY_5450_out0;
wire v$CARRY_5451_out0;
wire v$CARRY_5452_out0;
wire v$CARRY_5453_out0;
wire v$CARRY_5454_out0;
wire v$CARRY_5455_out0;
wire v$CARRY_5456_out0;
wire v$CARRY_5457_out0;
wire v$CARRY_5458_out0;
wire v$CARRY_5459_out0;
wire v$CARRY_5460_out0;
wire v$CARRY_5461_out0;
wire v$CARRY_5462_out0;
wire v$CARRY_5463_out0;
wire v$CARRY_5464_out0;
wire v$CARRY_5465_out0;
wire v$CARRY_5466_out0;
wire v$CARRY_5467_out0;
wire v$CARRY_5468_out0;
wire v$CARRY_5469_out0;
wire v$CARRY_5470_out0;
wire v$CARRY_5471_out0;
wire v$CARRY_5472_out0;
wire v$CARRY_5473_out0;
wire v$CARRY_5474_out0;
wire v$CARRY_5475_out0;
wire v$CARRY_5476_out0;
wire v$CARRY_5477_out0;
wire v$CARRY_5478_out0;
wire v$CARRY_5479_out0;
wire v$CARRY_5480_out0;
wire v$CARRY_5481_out0;
wire v$CARRY_5482_out0;
wire v$CARRY_5483_out0;
wire v$CARRY_5484_out0;
wire v$CARRY_5485_out0;
wire v$CARRY_5486_out0;
wire v$CARRY_5487_out0;
wire v$CARRY_5488_out0;
wire v$CARRY_5489_out0;
wire v$CARRY_5490_out0;
wire v$CARRY_5491_out0;
wire v$CARRY_5492_out0;
wire v$CARRY_5493_out0;
wire v$CARRY_5494_out0;
wire v$CARRY_5495_out0;
wire v$CARRY_5496_out0;
wire v$CARRY_5497_out0;
wire v$CARRY_5498_out0;
wire v$CARRY_5499_out0;
wire v$CARRY_5500_out0;
wire v$CARRY_5501_out0;
wire v$CARRY_5502_out0;
wire v$CARRY_5503_out0;
wire v$CARRY_5504_out0;
wire v$CARRY_5505_out0;
wire v$CARRY_5506_out0;
wire v$CARRY_5507_out0;
wire v$CARRY_5508_out0;
wire v$CARRY_5509_out0;
wire v$CARRY_5510_out0;
wire v$CARRY_5511_out0;
wire v$CARRY_5512_out0;
wire v$CARRY_5513_out0;
wire v$CARRY_5514_out0;
wire v$CARRY_5515_out0;
wire v$CARRY_5516_out0;
wire v$CARRY_5517_out0;
wire v$CARRY_5518_out0;
wire v$CARRY_5519_out0;
wire v$CARRY_5520_out0;
wire v$CARRY_5521_out0;
wire v$CARRY_5522_out0;
wire v$CARRY_5523_out0;
wire v$CARRY_5524_out0;
wire v$CARRY_5525_out0;
wire v$CARRY_5526_out0;
wire v$CARRY_5527_out0;
wire v$CARRY_5528_out0;
wire v$CARRY_5529_out0;
wire v$CARRY_5530_out0;
wire v$CARRY_5531_out0;
wire v$CARRY_5532_out0;
wire v$CARRY_5533_out0;
wire v$CARRY_5534_out0;
wire v$CARRY_5535_out0;
wire v$CARRY_5536_out0;
wire v$CARRY_5537_out0;
wire v$CARRY_5538_out0;
wire v$CARRY_5539_out0;
wire v$CARRY_5540_out0;
wire v$CARRY_5541_out0;
wire v$CARRY_5542_out0;
wire v$CARRY_5543_out0;
wire v$CARRY_5544_out0;
wire v$CARRY_5545_out0;
wire v$CARRY_5546_out0;
wire v$CARRY_5547_out0;
wire v$CARRY_5548_out0;
wire v$CARRY_5549_out0;
wire v$CARRY_5550_out0;
wire v$CARRY_5551_out0;
wire v$CARRY_5552_out0;
wire v$CARRY_5553_out0;
wire v$CARRY_5554_out0;
wire v$CARRY_5555_out0;
wire v$CARRY_5556_out0;
wire v$CARRY_5557_out0;
wire v$CARRY_5558_out0;
wire v$CARRY_5559_out0;
wire v$CARRY_5560_out0;
wire v$CARRY_5561_out0;
wire v$CARRY_5562_out0;
wire v$CARRY_5563_out0;
wire v$CARRY_5564_out0;
wire v$CARRY_5565_out0;
wire v$CARRY_5566_out0;
wire v$CARRY_5567_out0;
wire v$CARRY_5568_out0;
wire v$CARRY_5569_out0;
wire v$CARRY_5570_out0;
wire v$CARRY_5571_out0;
wire v$CARRY_5572_out0;
wire v$CARRY_5573_out0;
wire v$CARRY_5574_out0;
wire v$CARRY_5575_out0;
wire v$CARRY_5576_out0;
wire v$CARRY_5577_out0;
wire v$CARRY_5578_out0;
wire v$CARRY_5579_out0;
wire v$CARRY_5580_out0;
wire v$CARRY_5581_out0;
wire v$CARRY_5582_out0;
wire v$CARRY_5583_out0;
wire v$CARRY_5584_out0;
wire v$CARRY_5585_out0;
wire v$CARRY_5586_out0;
wire v$CARRY_5587_out0;
wire v$CARRY_5588_out0;
wire v$CARRY_5589_out0;
wire v$CARRY_5590_out0;
wire v$CARRY_5591_out0;
wire v$CARRY_5592_out0;
wire v$CARRY_5593_out0;
wire v$CARRY_5594_out0;
wire v$CARRY_5595_out0;
wire v$CARRY_5596_out0;
wire v$CARRY_5597_out0;
wire v$CARRY_5598_out0;
wire v$CARRY_5599_out0;
wire v$CARRY_5600_out0;
wire v$CARRY_5601_out0;
wire v$CARRY_5602_out0;
wire v$CARRY_5603_out0;
wire v$CARRY_5604_out0;
wire v$CARRY_5605_out0;
wire v$CARRY_5606_out0;
wire v$CARRY_5607_out0;
wire v$CARRY_5608_out0;
wire v$CARRY_5609_out0;
wire v$CARRY_5610_out0;
wire v$CARRY_5611_out0;
wire v$CARRY_5612_out0;
wire v$CARRY_5613_out0;
wire v$CARRY_5614_out0;
wire v$CARRY_5615_out0;
wire v$CARRY_5616_out0;
wire v$CARRY_5617_out0;
wire v$CARRY_5618_out0;
wire v$CARRY_5619_out0;
wire v$CARRY_5620_out0;
wire v$CARRY_5621_out0;
wire v$CARRY_5622_out0;
wire v$CARRY_5623_out0;
wire v$CARRY_5624_out0;
wire v$CARRY_5625_out0;
wire v$CARRY_5626_out0;
wire v$CARRY_5627_out0;
wire v$CARRY_5628_out0;
wire v$CARRY_5629_out0;
wire v$CARRY_5630_out0;
wire v$CARRY_5631_out0;
wire v$CARRY_5632_out0;
wire v$CARRY_5633_out0;
wire v$CARRY_5634_out0;
wire v$CARRY_5635_out0;
wire v$CARRY_5636_out0;
wire v$CARRY_5637_out0;
wire v$CARRY_5638_out0;
wire v$CARRY_5639_out0;
wire v$CARRY_5640_out0;
wire v$CARRY_5641_out0;
wire v$CARRY_5642_out0;
wire v$CARRY_5643_out0;
wire v$CARRY_5644_out0;
wire v$CARRY_5645_out0;
wire v$CARRY_5646_out0;
wire v$CARRY_5647_out0;
wire v$CARRY_5648_out0;
wire v$CARRY_5649_out0;
wire v$CARRY_5650_out0;
wire v$CARRY_5651_out0;
wire v$CARRY_5652_out0;
wire v$CARRY_5653_out0;
wire v$CARRY_5654_out0;
wire v$CARRY_5655_out0;
wire v$CARRY_5656_out0;
wire v$CARRY_5657_out0;
wire v$CARRY_5658_out0;
wire v$CARRY_5659_out0;
wire v$CARRY_5660_out0;
wire v$CARRY_5661_out0;
wire v$CARRY_5662_out0;
wire v$CARRY_5663_out0;
wire v$CARRY_5664_out0;
wire v$CARRY_5665_out0;
wire v$CARRY_5666_out0;
wire v$CARRY_5667_out0;
wire v$CARRY_5668_out0;
wire v$CARRY_5669_out0;
wire v$CARRY_5670_out0;
wire v$CARRY_5671_out0;
wire v$CARRY_5672_out0;
wire v$CARRY_5673_out0;
wire v$CARRY_5674_out0;
wire v$CARRY_5675_out0;
wire v$CARRY_5676_out0;
wire v$CARRY_5677_out0;
wire v$CARRY_5678_out0;
wire v$CARRY_5679_out0;
wire v$CARRY_5680_out0;
wire v$CARRY_5681_out0;
wire v$CARRY_5682_out0;
wire v$CARRY_5683_out0;
wire v$CARRY_5684_out0;
wire v$CARRY_5685_out0;
wire v$CARRY_5686_out0;
wire v$CARRY_5687_out0;
wire v$CARRY_5688_out0;
wire v$CARRY_5689_out0;
wire v$CARRY_5690_out0;
wire v$CARRY_5691_out0;
wire v$CARRY_5692_out0;
wire v$CARRY_5693_out0;
wire v$CARRY_5694_out0;
wire v$CARRY_5695_out0;
wire v$CARRY_5696_out0;
wire v$CARRY_5697_out0;
wire v$CARRY_5698_out0;
wire v$CARRY_5699_out0;
wire v$CARRY_5700_out0;
wire v$CARRY_5701_out0;
wire v$CARRY_5702_out0;
wire v$CARRY_5703_out0;
wire v$CARRY_5704_out0;
wire v$CARRY_5705_out0;
wire v$CARRY_5706_out0;
wire v$CARRY_5707_out0;
wire v$CARRY_5708_out0;
wire v$CARRY_5709_out0;
wire v$CARRY_5710_out0;
wire v$CARRY_5711_out0;
wire v$CARRY_5712_out0;
wire v$CARRY_5713_out0;
wire v$CARRY_5714_out0;
wire v$CARRY_5715_out0;
wire v$CARRY_5716_out0;
wire v$CARRY_5717_out0;
wire v$CARRY_5718_out0;
wire v$CARRY_5719_out0;
wire v$CARRY_5720_out0;
wire v$CARRY_5721_out0;
wire v$CARRY_5722_out0;
wire v$CARRY_5723_out0;
wire v$CARRY_5724_out0;
wire v$CARRY_5725_out0;
wire v$CARRY_5726_out0;
wire v$CARRY_5727_out0;
wire v$CARRY_5728_out0;
wire v$CARRY_5729_out0;
wire v$CARRY_5730_out0;
wire v$CARRY_5731_out0;
wire v$CARRY_5732_out0;
wire v$CARRY_5733_out0;
wire v$CARRY_5734_out0;
wire v$CARRY_5735_out0;
wire v$CARRY_5736_out0;
wire v$CARRY_5737_out0;
wire v$CARRY_5738_out0;
wire v$CARRY_5739_out0;
wire v$CARRY_5740_out0;
wire v$CARRY_5741_out0;
wire v$CARRY_5742_out0;
wire v$CARRY_5743_out0;
wire v$CARRY_5744_out0;
wire v$CARRY_5745_out0;
wire v$CARRY_5746_out0;
wire v$CARRY_5747_out0;
wire v$CARRY_5748_out0;
wire v$CARRY_5749_out0;
wire v$CARRY_5750_out0;
wire v$CARRY_5751_out0;
wire v$CARRY_5752_out0;
wire v$CARRY_5753_out0;
wire v$CARRY_5754_out0;
wire v$CARRY_5755_out0;
wire v$CARRY_5756_out0;
wire v$CARRY_5757_out0;
wire v$CARRY_5758_out0;
wire v$CARRY_5759_out0;
wire v$CARRY_5760_out0;
wire v$CARRY_5761_out0;
wire v$CARRY_5762_out0;
wire v$CARRY_5763_out0;
wire v$CARRY_5764_out0;
wire v$CARRY_5765_out0;
wire v$CARRY_5766_out0;
wire v$CARRY_5767_out0;
wire v$CARRY_5768_out0;
wire v$CARRY_5769_out0;
wire v$CARRY_5770_out0;
wire v$CARRY_5771_out0;
wire v$CARRY_5772_out0;
wire v$CARRY_5773_out0;
wire v$CARRY_5774_out0;
wire v$CARRY_5775_out0;
wire v$CARRY_5776_out0;
wire v$CARRY_5777_out0;
wire v$CARRY_5778_out0;
wire v$CARRY_5779_out0;
wire v$CARRY_5780_out0;
wire v$CARRY_5781_out0;
wire v$CARRY_5782_out0;
wire v$CARRY_5783_out0;
wire v$CARRY_5784_out0;
wire v$CARRY_5785_out0;
wire v$CARRY_5786_out0;
wire v$CARRY_5787_out0;
wire v$CARRY_5788_out0;
wire v$CARRY_5789_out0;
wire v$CIN_10000_out0;
wire v$CIN_10001_out0;
wire v$CIN_10002_out0;
wire v$CIN_10003_out0;
wire v$CIN_10004_out0;
wire v$CIN_10005_out0;
wire v$CIN_10006_out0;
wire v$CIN_10007_out0;
wire v$CIN_10008_out0;
wire v$CIN_10009_out0;
wire v$CIN_10010_out0;
wire v$CIN_10011_out0;
wire v$CIN_10012_out0;
wire v$CIN_10013_out0;
wire v$CIN_10014_out0;
wire v$CIN_10015_out0;
wire v$CIN_10016_out0;
wire v$CIN_10017_out0;
wire v$CIN_10018_out0;
wire v$CIN_10019_out0;
wire v$CIN_10020_out0;
wire v$CIN_10021_out0;
wire v$CIN_10022_out0;
wire v$CIN_10023_out0;
wire v$CIN_10024_out0;
wire v$CIN_10025_out0;
wire v$CIN_10026_out0;
wire v$CIN_10027_out0;
wire v$CIN_10028_out0;
wire v$CIN_10029_out0;
wire v$CIN_10030_out0;
wire v$CIN_10031_out0;
wire v$CIN_10032_out0;
wire v$CIN_10033_out0;
wire v$CIN_10034_out0;
wire v$CIN_10035_out0;
wire v$CIN_10036_out0;
wire v$CIN_10037_out0;
wire v$CIN_10038_out0;
wire v$CIN_10039_out0;
wire v$CIN_10040_out0;
wire v$CIN_10041_out0;
wire v$CIN_10042_out0;
wire v$CIN_10043_out0;
wire v$CIN_10044_out0;
wire v$CIN_10045_out0;
wire v$CIN_10046_out0;
wire v$CIN_10047_out0;
wire v$CIN_10048_out0;
wire v$CIN_10049_out0;
wire v$CIN_10050_out0;
wire v$CIN_10051_out0;
wire v$CIN_10052_out0;
wire v$CIN_10053_out0;
wire v$CIN_10054_out0;
wire v$CIN_10055_out0;
wire v$CIN_10056_out0;
wire v$CIN_10057_out0;
wire v$CIN_10058_out0;
wire v$CIN_10059_out0;
wire v$CIN_10060_out0;
wire v$CIN_10061_out0;
wire v$CIN_10062_out0;
wire v$CIN_10063_out0;
wire v$CIN_10064_out0;
wire v$CIN_10065_out0;
wire v$CIN_10066_out0;
wire v$CIN_10067_out0;
wire v$CIN_10068_out0;
wire v$CIN_10069_out0;
wire v$CIN_10070_out0;
wire v$CIN_10071_out0;
wire v$CIN_10072_out0;
wire v$CIN_10073_out0;
wire v$CIN_10074_out0;
wire v$CIN_10075_out0;
wire v$CIN_10076_out0;
wire v$CIN_10077_out0;
wire v$CIN_10078_out0;
wire v$CIN_10079_out0;
wire v$CIN_10080_out0;
wire v$CIN_10081_out0;
wire v$CIN_10082_out0;
wire v$CIN_10083_out0;
wire v$CIN_10084_out0;
wire v$CIN_10085_out0;
wire v$CIN_10086_out0;
wire v$CIN_10087_out0;
wire v$CIN_10088_out0;
wire v$CIN_10089_out0;
wire v$CIN_10090_out0;
wire v$CIN_10091_out0;
wire v$CIN_10092_out0;
wire v$CIN_10093_out0;
wire v$CIN_10094_out0;
wire v$CIN_10095_out0;
wire v$CIN_10096_out0;
wire v$CIN_10097_out0;
wire v$CIN_10098_out0;
wire v$CIN_10099_out0;
wire v$CIN_10100_out0;
wire v$CIN_10101_out0;
wire v$CIN_10102_out0;
wire v$CIN_10103_out0;
wire v$CIN_10104_out0;
wire v$CIN_10105_out0;
wire v$CIN_10106_out0;
wire v$CIN_10107_out0;
wire v$CIN_10108_out0;
wire v$CIN_10109_out0;
wire v$CIN_10110_out0;
wire v$CIN_10111_out0;
wire v$CIN_10112_out0;
wire v$CIN_10113_out0;
wire v$CIN_10114_out0;
wire v$CIN_10115_out0;
wire v$CIN_10116_out0;
wire v$CIN_10117_out0;
wire v$CIN_10118_out0;
wire v$CIN_10119_out0;
wire v$CIN_10120_out0;
wire v$CIN_10121_out0;
wire v$CIN_10122_out0;
wire v$CIN_10123_out0;
wire v$CIN_10124_out0;
wire v$CIN_10125_out0;
wire v$CIN_10126_out0;
wire v$CIN_10127_out0;
wire v$CIN_10128_out0;
wire v$CIN_10129_out0;
wire v$CIN_10130_out0;
wire v$CIN_10131_out0;
wire v$CIN_10132_out0;
wire v$CIN_10133_out0;
wire v$CIN_10134_out0;
wire v$CIN_10135_out0;
wire v$CIN_10136_out0;
wire v$CIN_10137_out0;
wire v$CIN_10138_out0;
wire v$CIN_10139_out0;
wire v$CIN_10140_out0;
wire v$CIN_10141_out0;
wire v$CIN_10142_out0;
wire v$CIN_10143_out0;
wire v$CIN_10144_out0;
wire v$CIN_10145_out0;
wire v$CIN_10146_out0;
wire v$CIN_10147_out0;
wire v$CIN_10148_out0;
wire v$CIN_10149_out0;
wire v$CIN_10150_out0;
wire v$CIN_10151_out0;
wire v$CIN_10152_out0;
wire v$CIN_10153_out0;
wire v$CIN_10154_out0;
wire v$CIN_10155_out0;
wire v$CIN_10156_out0;
wire v$CIN_10157_out0;
wire v$CIN_10158_out0;
wire v$CIN_10159_out0;
wire v$CIN_10160_out0;
wire v$CIN_10161_out0;
wire v$CIN_10162_out0;
wire v$CIN_10163_out0;
wire v$CIN_10164_out0;
wire v$CIN_10165_out0;
wire v$CIN_10166_out0;
wire v$CIN_10167_out0;
wire v$CIN_10168_out0;
wire v$CIN_10169_out0;
wire v$CIN_10170_out0;
wire v$CIN_10171_out0;
wire v$CIN_10172_out0;
wire v$CIN_10173_out0;
wire v$CIN_10174_out0;
wire v$CIN_10175_out0;
wire v$CIN_10176_out0;
wire v$CIN_10177_out0;
wire v$CIN_10178_out0;
wire v$CIN_10179_out0;
wire v$CIN_10180_out0;
wire v$CIN_10181_out0;
wire v$CIN_10182_out0;
wire v$CIN_10183_out0;
wire v$CIN_10184_out0;
wire v$CIN_10185_out0;
wire v$CIN_10186_out0;
wire v$CIN_10187_out0;
wire v$CIN_10188_out0;
wire v$CIN_10189_out0;
wire v$CIN_10190_out0;
wire v$CIN_10191_out0;
wire v$CIN_10192_out0;
wire v$CIN_10193_out0;
wire v$CIN_10194_out0;
wire v$CIN_10195_out0;
wire v$CIN_10196_out0;
wire v$CIN_10197_out0;
wire v$CIN_10198_out0;
wire v$CIN_10199_out0;
wire v$CIN_10200_out0;
wire v$CIN_10201_out0;
wire v$CIN_10202_out0;
wire v$CIN_10203_out0;
wire v$CIN_10204_out0;
wire v$CIN_10205_out0;
wire v$CIN_10206_out0;
wire v$CIN_10207_out0;
wire v$CIN_10208_out0;
wire v$CIN_10209_out0;
wire v$CIN_10210_out0;
wire v$CIN_10211_out0;
wire v$CIN_10212_out0;
wire v$CIN_10213_out0;
wire v$CIN_10214_out0;
wire v$CIN_10215_out0;
wire v$CIN_10216_out0;
wire v$CIN_10217_out0;
wire v$CIN_10218_out0;
wire v$CIN_10219_out0;
wire v$CIN_10220_out0;
wire v$CIN_10221_out0;
wire v$CIN_10222_out0;
wire v$CIN_10223_out0;
wire v$CIN_10224_out0;
wire v$CIN_10225_out0;
wire v$CIN_10226_out0;
wire v$CIN_10227_out0;
wire v$CIN_10228_out0;
wire v$CIN_10229_out0;
wire v$CIN_10230_out0;
wire v$CIN_10231_out0;
wire v$CIN_10232_out0;
wire v$CIN_10233_out0;
wire v$CIN_10234_out0;
wire v$CIN_10235_out0;
wire v$CIN_10236_out0;
wire v$CIN_10237_out0;
wire v$CIN_10238_out0;
wire v$CIN_10239_out0;
wire v$CIN_10240_out0;
wire v$CIN_10241_out0;
wire v$CIN_10242_out0;
wire v$CIN_10243_out0;
wire v$CIN_10244_out0;
wire v$CIN_10245_out0;
wire v$CIN_10246_out0;
wire v$CIN_10247_out0;
wire v$CIN_10248_out0;
wire v$CIN_10249_out0;
wire v$CIN_10250_out0;
wire v$CIN_10251_out0;
wire v$CIN_10252_out0;
wire v$CIN_10253_out0;
wire v$CIN_10254_out0;
wire v$CIN_10255_out0;
wire v$CIN_9808_out0;
wire v$CIN_9809_out0;
wire v$CIN_9810_out0;
wire v$CIN_9811_out0;
wire v$CIN_9812_out0;
wire v$CIN_9813_out0;
wire v$CIN_9814_out0;
wire v$CIN_9815_out0;
wire v$CIN_9816_out0;
wire v$CIN_9817_out0;
wire v$CIN_9818_out0;
wire v$CIN_9819_out0;
wire v$CIN_9820_out0;
wire v$CIN_9821_out0;
wire v$CIN_9822_out0;
wire v$CIN_9823_out0;
wire v$CIN_9824_out0;
wire v$CIN_9825_out0;
wire v$CIN_9826_out0;
wire v$CIN_9827_out0;
wire v$CIN_9828_out0;
wire v$CIN_9829_out0;
wire v$CIN_9830_out0;
wire v$CIN_9831_out0;
wire v$CIN_9832_out0;
wire v$CIN_9833_out0;
wire v$CIN_9834_out0;
wire v$CIN_9835_out0;
wire v$CIN_9836_out0;
wire v$CIN_9837_out0;
wire v$CIN_9838_out0;
wire v$CIN_9839_out0;
wire v$CIN_9840_out0;
wire v$CIN_9841_out0;
wire v$CIN_9842_out0;
wire v$CIN_9843_out0;
wire v$CIN_9844_out0;
wire v$CIN_9845_out0;
wire v$CIN_9846_out0;
wire v$CIN_9847_out0;
wire v$CIN_9848_out0;
wire v$CIN_9849_out0;
wire v$CIN_9850_out0;
wire v$CIN_9851_out0;
wire v$CIN_9852_out0;
wire v$CIN_9853_out0;
wire v$CIN_9854_out0;
wire v$CIN_9855_out0;
wire v$CIN_9856_out0;
wire v$CIN_9857_out0;
wire v$CIN_9858_out0;
wire v$CIN_9859_out0;
wire v$CIN_9860_out0;
wire v$CIN_9861_out0;
wire v$CIN_9862_out0;
wire v$CIN_9863_out0;
wire v$CIN_9864_out0;
wire v$CIN_9865_out0;
wire v$CIN_9866_out0;
wire v$CIN_9867_out0;
wire v$CIN_9868_out0;
wire v$CIN_9869_out0;
wire v$CIN_9870_out0;
wire v$CIN_9871_out0;
wire v$CIN_9872_out0;
wire v$CIN_9873_out0;
wire v$CIN_9874_out0;
wire v$CIN_9875_out0;
wire v$CIN_9876_out0;
wire v$CIN_9877_out0;
wire v$CIN_9878_out0;
wire v$CIN_9879_out0;
wire v$CIN_9880_out0;
wire v$CIN_9881_out0;
wire v$CIN_9882_out0;
wire v$CIN_9883_out0;
wire v$CIN_9884_out0;
wire v$CIN_9885_out0;
wire v$CIN_9886_out0;
wire v$CIN_9887_out0;
wire v$CIN_9888_out0;
wire v$CIN_9889_out0;
wire v$CIN_9890_out0;
wire v$CIN_9891_out0;
wire v$CIN_9892_out0;
wire v$CIN_9893_out0;
wire v$CIN_9894_out0;
wire v$CIN_9895_out0;
wire v$CIN_9896_out0;
wire v$CIN_9897_out0;
wire v$CIN_9898_out0;
wire v$CIN_9899_out0;
wire v$CIN_9900_out0;
wire v$CIN_9901_out0;
wire v$CIN_9902_out0;
wire v$CIN_9903_out0;
wire v$CIN_9904_out0;
wire v$CIN_9905_out0;
wire v$CIN_9906_out0;
wire v$CIN_9907_out0;
wire v$CIN_9908_out0;
wire v$CIN_9909_out0;
wire v$CIN_9910_out0;
wire v$CIN_9911_out0;
wire v$CIN_9912_out0;
wire v$CIN_9913_out0;
wire v$CIN_9914_out0;
wire v$CIN_9915_out0;
wire v$CIN_9916_out0;
wire v$CIN_9917_out0;
wire v$CIN_9918_out0;
wire v$CIN_9919_out0;
wire v$CIN_9920_out0;
wire v$CIN_9921_out0;
wire v$CIN_9922_out0;
wire v$CIN_9923_out0;
wire v$CIN_9924_out0;
wire v$CIN_9925_out0;
wire v$CIN_9926_out0;
wire v$CIN_9927_out0;
wire v$CIN_9928_out0;
wire v$CIN_9929_out0;
wire v$CIN_9930_out0;
wire v$CIN_9931_out0;
wire v$CIN_9932_out0;
wire v$CIN_9933_out0;
wire v$CIN_9934_out0;
wire v$CIN_9935_out0;
wire v$CIN_9936_out0;
wire v$CIN_9937_out0;
wire v$CIN_9938_out0;
wire v$CIN_9939_out0;
wire v$CIN_9940_out0;
wire v$CIN_9941_out0;
wire v$CIN_9942_out0;
wire v$CIN_9943_out0;
wire v$CIN_9944_out0;
wire v$CIN_9945_out0;
wire v$CIN_9946_out0;
wire v$CIN_9947_out0;
wire v$CIN_9948_out0;
wire v$CIN_9949_out0;
wire v$CIN_9950_out0;
wire v$CIN_9951_out0;
wire v$CIN_9952_out0;
wire v$CIN_9953_out0;
wire v$CIN_9954_out0;
wire v$CIN_9955_out0;
wire v$CIN_9956_out0;
wire v$CIN_9957_out0;
wire v$CIN_9958_out0;
wire v$CIN_9959_out0;
wire v$CIN_9960_out0;
wire v$CIN_9961_out0;
wire v$CIN_9962_out0;
wire v$CIN_9963_out0;
wire v$CIN_9964_out0;
wire v$CIN_9965_out0;
wire v$CIN_9966_out0;
wire v$CIN_9967_out0;
wire v$CIN_9968_out0;
wire v$CIN_9969_out0;
wire v$CIN_9970_out0;
wire v$CIN_9971_out0;
wire v$CIN_9972_out0;
wire v$CIN_9973_out0;
wire v$CIN_9974_out0;
wire v$CIN_9975_out0;
wire v$CIN_9976_out0;
wire v$CIN_9977_out0;
wire v$CIN_9978_out0;
wire v$CIN_9979_out0;
wire v$CIN_9980_out0;
wire v$CIN_9981_out0;
wire v$CIN_9982_out0;
wire v$CIN_9983_out0;
wire v$CIN_9984_out0;
wire v$CIN_9985_out0;
wire v$CIN_9986_out0;
wire v$CIN_9987_out0;
wire v$CIN_9988_out0;
wire v$CIN_9989_out0;
wire v$CIN_9990_out0;
wire v$CIN_9991_out0;
wire v$CIN_9992_out0;
wire v$CIN_9993_out0;
wire v$CIN_9994_out0;
wire v$CIN_9995_out0;
wire v$CIN_9996_out0;
wire v$CIN_9997_out0;
wire v$CIN_9998_out0;
wire v$CIN_9999_out0;
wire v$CMP_13609_out0;
wire v$CMP_13610_out0;
wire v$CMP_3805_out0;
wire v$CMP_3806_out0;
wire v$CMP_8646_out0;
wire v$CMP_8647_out0;
wire v$COUT_1000_out0;
wire v$COUT_1001_out0;
wire v$COUT_1002_out0;
wire v$COUT_1003_out0;
wire v$COUT_1004_out0;
wire v$COUT_1005_out0;
wire v$COUT_1006_out0;
wire v$COUT_1007_out0;
wire v$COUT_1008_out0;
wire v$COUT_1009_out0;
wire v$COUT_1010_out0;
wire v$COUT_1011_out0;
wire v$COUT_1012_out0;
wire v$COUT_1013_out0;
wire v$COUT_1014_out0;
wire v$COUT_1015_out0;
wire v$COUT_1016_out0;
wire v$COUT_1017_out0;
wire v$COUT_1018_out0;
wire v$COUT_1019_out0;
wire v$COUT_1020_out0;
wire v$COUT_1021_out0;
wire v$COUT_1022_out0;
wire v$COUT_1023_out0;
wire v$COUT_1024_out0;
wire v$COUT_1025_out0;
wire v$COUT_1026_out0;
wire v$COUT_1027_out0;
wire v$COUT_1028_out0;
wire v$COUT_1029_out0;
wire v$COUT_1030_out0;
wire v$COUT_1031_out0;
wire v$COUT_1032_out0;
wire v$COUT_1033_out0;
wire v$COUT_1034_out0;
wire v$COUT_1035_out0;
wire v$COUT_1036_out0;
wire v$COUT_1037_out0;
wire v$COUT_1038_out0;
wire v$COUT_1039_out0;
wire v$COUT_1040_out0;
wire v$COUT_1041_out0;
wire v$COUT_1042_out0;
wire v$COUT_1043_out0;
wire v$COUT_1044_out0;
wire v$COUT_1045_out0;
wire v$COUT_1046_out0;
wire v$COUT_1047_out0;
wire v$COUT_1048_out0;
wire v$COUT_1049_out0;
wire v$COUT_1050_out0;
wire v$COUT_1051_out0;
wire v$COUT_1052_out0;
wire v$COUT_1053_out0;
wire v$COUT_10547_out0;
wire v$COUT_10548_out0;
wire v$COUT_1054_out0;
wire v$COUT_1055_out0;
wire v$COUT_1056_out0;
wire v$COUT_1057_out0;
wire v$COUT_1058_out0;
wire v$COUT_1059_out0;
wire v$COUT_1060_out0;
wire v$COUT_1061_out0;
wire v$COUT_1062_out0;
wire v$COUT_1063_out0;
wire v$COUT_1064_out0;
wire v$COUT_1065_out0;
wire v$COUT_1066_out0;
wire v$COUT_1067_out0;
wire v$COUT_1068_out0;
wire v$COUT_1069_out0;
wire v$COUT_1070_out0;
wire v$COUT_1071_out0;
wire v$COUT_1072_out0;
wire v$COUT_1073_out0;
wire v$COUT_1074_out0;
wire v$COUT_1075_out0;
wire v$COUT_1076_out0;
wire v$COUT_1077_out0;
wire v$COUT_1078_out0;
wire v$COUT_1079_out0;
wire v$COUT_1080_out0;
wire v$COUT_1081_out0;
wire v$COUT_1082_out0;
wire v$COUT_1083_out0;
wire v$COUT_1084_out0;
wire v$COUT_1085_out0;
wire v$COUT_1086_out0;
wire v$COUT_1087_out0;
wire v$COUT_1088_out0;
wire v$COUT_1089_out0;
wire v$COUT_1090_out0;
wire v$COUT_1091_out0;
wire v$COUT_1092_out0;
wire v$COUT_1093_out0;
wire v$COUT_1094_out0;
wire v$COUT_1095_out0;
wire v$COUT_1096_out0;
wire v$COUT_1097_out0;
wire v$COUT_1098_out0;
wire v$COUT_1099_out0;
wire v$COUT_1100_out0;
wire v$COUT_1101_out0;
wire v$COUT_1102_out0;
wire v$COUT_1103_out0;
wire v$COUT_1104_out0;
wire v$COUT_1105_out0;
wire v$COUT_1106_out0;
wire v$COUT_1107_out0;
wire v$COUT_1108_out0;
wire v$COUT_1109_out0;
wire v$COUT_1110_out0;
wire v$COUT_1111_out0;
wire v$COUT_1112_out0;
wire v$COUT_1113_out0;
wire v$COUT_1114_out0;
wire v$COUT_1115_out0;
wire v$COUT_1116_out0;
wire v$COUT_1117_out0;
wire v$COUT_1118_out0;
wire v$COUT_1119_out0;
wire v$COUT_1120_out0;
wire v$COUT_1121_out0;
wire v$COUT_1122_out0;
wire v$COUT_1123_out0;
wire v$COUT_1124_out0;
wire v$COUT_1125_out0;
wire v$COUT_1126_out0;
wire v$COUT_1127_out0;
wire v$COUT_1128_out0;
wire v$COUT_1129_out0;
wire v$COUT_1130_out0;
wire v$COUT_1131_out0;
wire v$COUT_1132_out0;
wire v$COUT_1133_out0;
wire v$COUT_1134_out0;
wire v$COUT_2725_out0;
wire v$COUT_3895_out0;
wire v$COUT_3896_out0;
wire v$COUT_687_out0;
wire v$COUT_688_out0;
wire v$COUT_689_out0;
wire v$COUT_690_out0;
wire v$COUT_691_out0;
wire v$COUT_692_out0;
wire v$COUT_693_out0;
wire v$COUT_694_out0;
wire v$COUT_695_out0;
wire v$COUT_696_out0;
wire v$COUT_697_out0;
wire v$COUT_698_out0;
wire v$COUT_699_out0;
wire v$COUT_700_out0;
wire v$COUT_701_out0;
wire v$COUT_702_out0;
wire v$COUT_703_out0;
wire v$COUT_704_out0;
wire v$COUT_705_out0;
wire v$COUT_706_out0;
wire v$COUT_707_out0;
wire v$COUT_708_out0;
wire v$COUT_709_out0;
wire v$COUT_70_out0;
wire v$COUT_710_out0;
wire v$COUT_711_out0;
wire v$COUT_712_out0;
wire v$COUT_713_out0;
wire v$COUT_714_out0;
wire v$COUT_715_out0;
wire v$COUT_716_out0;
wire v$COUT_717_out0;
wire v$COUT_718_out0;
wire v$COUT_719_out0;
wire v$COUT_71_out0;
wire v$COUT_720_out0;
wire v$COUT_721_out0;
wire v$COUT_722_out0;
wire v$COUT_723_out0;
wire v$COUT_724_out0;
wire v$COUT_725_out0;
wire v$COUT_726_out0;
wire v$COUT_727_out0;
wire v$COUT_728_out0;
wire v$COUT_729_out0;
wire v$COUT_730_out0;
wire v$COUT_731_out0;
wire v$COUT_732_out0;
wire v$COUT_733_out0;
wire v$COUT_734_out0;
wire v$COUT_735_out0;
wire v$COUT_736_out0;
wire v$COUT_737_out0;
wire v$COUT_738_out0;
wire v$COUT_739_out0;
wire v$COUT_740_out0;
wire v$COUT_741_out0;
wire v$COUT_742_out0;
wire v$COUT_743_out0;
wire v$COUT_744_out0;
wire v$COUT_745_out0;
wire v$COUT_746_out0;
wire v$COUT_747_out0;
wire v$COUT_748_out0;
wire v$COUT_749_out0;
wire v$COUT_750_out0;
wire v$COUT_751_out0;
wire v$COUT_752_out0;
wire v$COUT_753_out0;
wire v$COUT_754_out0;
wire v$COUT_755_out0;
wire v$COUT_756_out0;
wire v$COUT_757_out0;
wire v$COUT_758_out0;
wire v$COUT_759_out0;
wire v$COUT_760_out0;
wire v$COUT_761_out0;
wire v$COUT_762_out0;
wire v$COUT_763_out0;
wire v$COUT_764_out0;
wire v$COUT_765_out0;
wire v$COUT_766_out0;
wire v$COUT_767_out0;
wire v$COUT_768_out0;
wire v$COUT_769_out0;
wire v$COUT_770_out0;
wire v$COUT_771_out0;
wire v$COUT_772_out0;
wire v$COUT_773_out0;
wire v$COUT_774_out0;
wire v$COUT_775_out0;
wire v$COUT_776_out0;
wire v$COUT_777_out0;
wire v$COUT_778_out0;
wire v$COUT_779_out0;
wire v$COUT_780_out0;
wire v$COUT_781_out0;
wire v$COUT_782_out0;
wire v$COUT_783_out0;
wire v$COUT_784_out0;
wire v$COUT_785_out0;
wire v$COUT_786_out0;
wire v$COUT_787_out0;
wire v$COUT_788_out0;
wire v$COUT_789_out0;
wire v$COUT_790_out0;
wire v$COUT_791_out0;
wire v$COUT_792_out0;
wire v$COUT_793_out0;
wire v$COUT_794_out0;
wire v$COUT_795_out0;
wire v$COUT_796_out0;
wire v$COUT_797_out0;
wire v$COUT_798_out0;
wire v$COUT_799_out0;
wire v$COUT_800_out0;
wire v$COUT_801_out0;
wire v$COUT_802_out0;
wire v$COUT_803_out0;
wire v$COUT_804_out0;
wire v$COUT_805_out0;
wire v$COUT_806_out0;
wire v$COUT_807_out0;
wire v$COUT_808_out0;
wire v$COUT_809_out0;
wire v$COUT_810_out0;
wire v$COUT_811_out0;
wire v$COUT_812_out0;
wire v$COUT_813_out0;
wire v$COUT_814_out0;
wire v$COUT_815_out0;
wire v$COUT_816_out0;
wire v$COUT_817_out0;
wire v$COUT_818_out0;
wire v$COUT_819_out0;
wire v$COUT_820_out0;
wire v$COUT_821_out0;
wire v$COUT_822_out0;
wire v$COUT_823_out0;
wire v$COUT_824_out0;
wire v$COUT_825_out0;
wire v$COUT_826_out0;
wire v$COUT_827_out0;
wire v$COUT_828_out0;
wire v$COUT_829_out0;
wire v$COUT_830_out0;
wire v$COUT_831_out0;
wire v$COUT_832_out0;
wire v$COUT_833_out0;
wire v$COUT_834_out0;
wire v$COUT_835_out0;
wire v$COUT_836_out0;
wire v$COUT_837_out0;
wire v$COUT_838_out0;
wire v$COUT_839_out0;
wire v$COUT_840_out0;
wire v$COUT_841_out0;
wire v$COUT_842_out0;
wire v$COUT_843_out0;
wire v$COUT_844_out0;
wire v$COUT_845_out0;
wire v$COUT_846_out0;
wire v$COUT_847_out0;
wire v$COUT_848_out0;
wire v$COUT_849_out0;
wire v$COUT_850_out0;
wire v$COUT_851_out0;
wire v$COUT_852_out0;
wire v$COUT_853_out0;
wire v$COUT_854_out0;
wire v$COUT_855_out0;
wire v$COUT_856_out0;
wire v$COUT_857_out0;
wire v$COUT_858_out0;
wire v$COUT_859_out0;
wire v$COUT_860_out0;
wire v$COUT_861_out0;
wire v$COUT_862_out0;
wire v$COUT_863_out0;
wire v$COUT_864_out0;
wire v$COUT_865_out0;
wire v$COUT_866_out0;
wire v$COUT_867_out0;
wire v$COUT_868_out0;
wire v$COUT_869_out0;
wire v$COUT_870_out0;
wire v$COUT_871_out0;
wire v$COUT_872_out0;
wire v$COUT_873_out0;
wire v$COUT_874_out0;
wire v$COUT_875_out0;
wire v$COUT_876_out0;
wire v$COUT_877_out0;
wire v$COUT_878_out0;
wire v$COUT_879_out0;
wire v$COUT_880_out0;
wire v$COUT_881_out0;
wire v$COUT_882_out0;
wire v$COUT_883_out0;
wire v$COUT_884_out0;
wire v$COUT_885_out0;
wire v$COUT_886_out0;
wire v$COUT_887_out0;
wire v$COUT_888_out0;
wire v$COUT_889_out0;
wire v$COUT_890_out0;
wire v$COUT_891_out0;
wire v$COUT_892_out0;
wire v$COUT_893_out0;
wire v$COUT_894_out0;
wire v$COUT_895_out0;
wire v$COUT_896_out0;
wire v$COUT_897_out0;
wire v$COUT_898_out0;
wire v$COUT_899_out0;
wire v$COUT_900_out0;
wire v$COUT_901_out0;
wire v$COUT_902_out0;
wire v$COUT_903_out0;
wire v$COUT_904_out0;
wire v$COUT_905_out0;
wire v$COUT_906_out0;
wire v$COUT_907_out0;
wire v$COUT_908_out0;
wire v$COUT_909_out0;
wire v$COUT_910_out0;
wire v$COUT_911_out0;
wire v$COUT_912_out0;
wire v$COUT_913_out0;
wire v$COUT_914_out0;
wire v$COUT_915_out0;
wire v$COUT_916_out0;
wire v$COUT_917_out0;
wire v$COUT_918_out0;
wire v$COUT_919_out0;
wire v$COUT_920_out0;
wire v$COUT_921_out0;
wire v$COUT_922_out0;
wire v$COUT_923_out0;
wire v$COUT_924_out0;
wire v$COUT_925_out0;
wire v$COUT_926_out0;
wire v$COUT_927_out0;
wire v$COUT_928_out0;
wire v$COUT_929_out0;
wire v$COUT_930_out0;
wire v$COUT_931_out0;
wire v$COUT_932_out0;
wire v$COUT_933_out0;
wire v$COUT_934_out0;
wire v$COUT_935_out0;
wire v$COUT_936_out0;
wire v$COUT_937_out0;
wire v$COUT_938_out0;
wire v$COUT_939_out0;
wire v$COUT_940_out0;
wire v$COUT_941_out0;
wire v$COUT_942_out0;
wire v$COUT_943_out0;
wire v$COUT_944_out0;
wire v$COUT_945_out0;
wire v$COUT_946_out0;
wire v$COUT_947_out0;
wire v$COUT_948_out0;
wire v$COUT_949_out0;
wire v$COUT_950_out0;
wire v$COUT_951_out0;
wire v$COUT_952_out0;
wire v$COUT_953_out0;
wire v$COUT_954_out0;
wire v$COUT_955_out0;
wire v$COUT_956_out0;
wire v$COUT_957_out0;
wire v$COUT_958_out0;
wire v$COUT_959_out0;
wire v$COUT_960_out0;
wire v$COUT_961_out0;
wire v$COUT_962_out0;
wire v$COUT_963_out0;
wire v$COUT_964_out0;
wire v$COUT_965_out0;
wire v$COUT_966_out0;
wire v$COUT_967_out0;
wire v$COUT_968_out0;
wire v$COUT_969_out0;
wire v$COUT_970_out0;
wire v$COUT_971_out0;
wire v$COUT_972_out0;
wire v$COUT_973_out0;
wire v$COUT_974_out0;
wire v$COUT_975_out0;
wire v$COUT_976_out0;
wire v$COUT_977_out0;
wire v$COUT_978_out0;
wire v$COUT_979_out0;
wire v$COUT_980_out0;
wire v$COUT_981_out0;
wire v$COUT_982_out0;
wire v$COUT_983_out0;
wire v$COUT_984_out0;
wire v$COUT_985_out0;
wire v$COUT_986_out0;
wire v$COUT_987_out0;
wire v$COUT_988_out0;
wire v$COUT_989_out0;
wire v$COUT_990_out0;
wire v$COUT_991_out0;
wire v$COUT_992_out0;
wire v$COUT_993_out0;
wire v$COUT_994_out0;
wire v$COUT_995_out0;
wire v$COUT_996_out0;
wire v$COUT_997_out0;
wire v$COUT_998_out0;
wire v$COUT_999_out0;
wire v$C_13767_out0;
wire v$C_13768_out0;
wire v$C_238_out0;
wire v$C_239_out0;
wire v$C_3197_out0;
wire v$C_3198_out0;
wire v$C_3207_out0;
wire v$C_3208_out0;
wire v$C_379_out0;
wire v$C_380_out0;
wire v$C_4848_out0;
wire v$C_4849_out0;
wire v$C_8648_out0;
wire v$C_8649_out0;
wire v$C_8653_out0;
wire v$C_8654_out0;
wire v$D1_8842_out0;
wire v$D1_8842_out1;
wire v$D1_8842_out2;
wire v$D1_8842_out3;
wire v$D1_8843_out0;
wire v$D1_8843_out1;
wire v$D1_8843_out2;
wire v$D1_8843_out3;
wire v$DIV$INSTRUCTION_11296_out0;
wire v$DIV$INSTRUCTION_11297_out0;
wire v$DIV$INSTRUCTION_13635_out0;
wire v$DIV$INSTRUCTION_13636_out0;
wire v$DIV$INSTRUCTION_3296_out0;
wire v$DIV$INSTRUCTION_3297_out0;
wire v$DIV$INSTRUCTION_4614_out0;
wire v$DIV$INSTRUCTION_4615_out0;
wire v$DIV$INST_2324_out0;
wire v$DIV$INST_2325_out0;
wire v$DONE$RECEIVING_3084_out0;
wire v$DONE$RECEIVING_5857_out0;
wire v$D_7679_out0;
wire v$D_7680_out0;
wire v$D_7681_out0;
wire v$D_7682_out0;
wire v$D_7683_out0;
wire v$D_7684_out0;
wire v$D_7685_out0;
wire v$D_7686_out0;
wire v$D_7687_out0;
wire v$D_7688_out0;
wire v$D_7689_out0;
wire v$D_7690_out0;
wire v$D_7691_out0;
wire v$D_7692_out0;
wire v$D_7693_out0;
wire v$D_7694_out0;
wire v$EN$STALL_10344_out0;
wire v$EN$STALL_13747_out0;
wire v$ENABLE_1757_out0;
wire v$ENABLE_2018_out0;
wire v$ENABLE_2019_out0;
wire v$ENABLE_2020_out0;
wire v$ENABLE_2021_out0;
wire v$ENABLE_2651_out0;
wire v$EN_10451_out0;
wire v$EN_10452_out0;
wire v$EN_10453_out0;
wire v$EN_10454_out0;
wire v$EN_10474_out0;
wire v$EN_10475_out0;
wire v$EN_13181_out0;
wire v$EN_13182_out0;
wire v$EN_2330_out0;
wire v$EN_2331_out0;
wire v$EN_2445_out0;
wire v$EN_2446_out0;
wire v$EN_2919_out0;
wire v$EN_2920_out0;
wire v$EN_2921_out0;
wire v$EN_2922_out0;
wire v$EN_2923_out0;
wire v$EN_2924_out0;
wire v$EN_2925_out0;
wire v$EN_2926_out0;
wire v$EN_2927_out0;
wire v$EN_2928_out0;
wire v$EN_2929_out0;
wire v$EN_2930_out0;
wire v$EN_2931_out0;
wire v$EN_2932_out0;
wire v$EN_2933_out0;
wire v$EN_2934_out0;
wire v$EN_4485_out0;
wire v$EN_4593_out0;
wire v$EN_4594_out0;
wire v$EN_7093_out0;
wire v$EN_7094_out0;
wire v$EQ01_10510_out0;
wire v$EQ01_10511_out0;
wire v$EQ10_2320_out0;
wire v$EQ10_2321_out0;
wire v$EQ11_2456_out0;
wire v$EQ11_2457_out0;
wire v$EQ11_4465_out0;
wire v$EQ11_4466_out0;
wire v$EQ1_10329_out0;
wire v$EQ1_1157_out0;
wire v$EQ1_1158_out0;
wire v$EQ1_13433_out0;
wire v$EQ1_13434_out0;
wire v$EQ1_1857_out0;
wire v$EQ1_1858_out0;
wire v$EQ1_2540_out0;
wire v$EQ1_2541_out0;
wire v$EQ1_2597_out0;
wire v$EQ1_2598_out0;
wire v$EQ1_2675_out0;
wire v$EQ1_2676_out0;
wire v$EQ1_315_out0;
wire v$EQ1_316_out0;
wire v$EQ1_3344_out0;
wire v$EQ1_6956_out0;
wire v$EQ1_6957_out0;
wire v$EQ1_7098_out0;
wire v$EQ1_7099_out0;
wire v$EQ2_10347_out0;
wire v$EQ2_10348_out0;
wire v$EQ2_10771_out0;
wire v$EQ2_10772_out0;
wire v$EQ2_10981_out0;
wire v$EQ2_11254_out0;
wire v$EQ2_11255_out0;
wire v$EQ2_1753_out0;
wire v$EQ2_1754_out0;
wire v$EQ2_7091_out0;
wire v$EQ2_7092_out0;
wire v$EQ2_8_out0;
wire v$EQ2_9795_out0;
wire v$EQ2_9_out0;
wire v$EQ3_11044_out0;
wire v$EQ3_11045_out0;
wire v$EQ3_13504_out0;
wire v$EQ3_13505_out0;
wire v$EQ3_2966_out0;
wire v$EQ3_2967_out0;
wire v$EQ3_5861_out0;
wire v$EQ3_7126_out0;
wire v$EQ3_7127_out0;
wire v$EQ3_7145_out0;
wire v$EQ3_7146_out0;
wire v$EQ4_10345_out0;
wire v$EQ4_10346_out0;
wire v$EQ4_1142_out0;
wire v$EQ4_2149_out0;
wire v$EQ4_3227_out0;
wire v$EQ4_3228_out0;
wire v$EQ4_611_out0;
wire v$EQ4_612_out0;
wire v$EQ5_10364_out0;
wire v$EQ5_10365_out0;
wire v$EQ5_4860_out0;
wire v$EQ5_4861_out0;
wire v$EQ6_1686_out0;
wire v$EQ6_1687_out0;
wire v$EQ6_1966_out0;
wire v$EQ6_1967_out0;
wire v$EQ6_19_out0;
wire v$EQ6_3257_out0;
wire v$EQ7_10399_out0;
wire v$EQ7_10400_out0;
wire v$EQ7_13769_out0;
wire v$EQ7_3307_out0;
wire v$EQ7_3308_out0;
wire v$EQ8_10804_out0;
wire v$EQ8_10805_out0;
wire v$EQ8_2453_out0;
wire v$EQ8_2454_out0;
wire v$EQ8_2874_out0;
wire v$EQ8_2951_out0;
wire v$EQ8_2952_out0;
wire v$EQ9_2007_out0;
wire v$EQ9_2390_out0;
wire v$EQ9_2391_out0;
wire v$EQ9_4842_out0;
wire v$EQ9_4843_out0;
wire v$EQ_100_out0;
wire v$EQ_101_out0;
wire v$EQ_2591_out0;
wire v$EQ_2592_out0;
wire v$EQ_3821_out0;
wire v$EQ_3822_out0;
wire v$EQ_4835_out0;
wire v$EQ_4836_out0;
wire v$EXEC10_2329_out0;
wire v$EXEC10_8812_out0;
wire v$EXEC11_2830_out0;
wire v$EXEC11_4528_out0;
wire v$EXEC1LS_10506_out0;
wire v$EXEC1LS_10507_out0;
wire v$EXEC1LS_10703_out0;
wire v$EXEC1LS_10704_out0;
wire v$EXEC1LS_10843_out0;
wire v$EXEC1LS_10844_out0;
wire v$EXEC1LS_430_out0;
wire v$EXEC1LS_431_out0;
wire v$EXEC1LS_4697_out0;
wire v$EXEC1LS_4698_out0;
wire v$EXEC1LS_6795_out0;
wire v$EXEC1LS_6796_out0;
wire v$EXEC1_10763_out0;
wire v$EXEC1_10764_out0;
wire v$EXEC1_1863_out0;
wire v$EXEC1_1864_out0;
wire v$EXEC1_20_out0;
wire v$EXEC1_21_out0;
wire v$EXEC1_2634_out0;
wire v$EXEC1_2635_out0;
wire v$EXEC1_3038_out0;
wire v$EXEC1_3039_out0;
wire v$EXEC1_7029_out0;
wire v$EXEC1_7030_out0;
wire v$EXEC1_7128_out0;
wire v$EXEC1_7129_out0;
wire v$EXEC20_629_out0;
wire v$EXEC2LS_10549_out0;
wire v$EXEC2LS_10979_out0;
wire v$EXEC2LS_10980_out0;
wire v$EXEC2LS_13558_out0;
wire v$EXEC2LS_13559_out0;
wire v$EXEC2LS_2844_out0;
wire v$EXEC2LS_2845_out0;
wire v$EXEC2LS_3081_out0;
wire v$EXEC2LS_3082_out0;
wire v$EXEC2LS_3188_out0;
wire v$EXEC2LS_3189_out0;
wire v$EXEC2LS_3231_out0;
wire v$EXEC2LS_3232_out0;
wire v$EXEC2_2010_out0;
wire v$EXEC2_2011_out0;
wire v$EXEC2_2110_out0;
wire v$EXEC2_2111_out0;
wire v$EXEC2_2647_out0;
wire v$EXEC2_2648_out0;
wire v$EXEC2_3170_out0;
wire v$EXEC2_3171_out0;
wire v$EXEC2_3241_out0;
wire v$EXEC2_3242_out0;
wire v$EXEC2_441_out0;
wire v$EXEC2_442_out0;
wire v$EXEC2_7181_out0;
wire v$EXEC2_7182_out0;
wire v$EXP1_13488_out0;
wire v$EXP1_13489_out0;
wire v$FLAOTING$INSTRUCTION_1859_out0;
wire v$FLAOTING$INSTRUCTION_1860_out0;
wire v$FLOAT$INST16_13443_out0;
wire v$FLOAT$INST16_13444_out0;
wire v$FLOAT$INST_2955_out0;
wire v$FLOAT$INST_2956_out0;
wire v$FLOATING$EN$ALU_634_out0;
wire v$FLOATING$EN$ALU_635_out0;
wire v$FLOATING$INSTRUCTION_10391_out0;
wire v$FLOATING$INSTRUCTION_10392_out0;
wire v$FLOATING$INS_13797_out0;
wire v$FLOATING$INS_13798_out0;
wire v$FLOAT_4603_out0;
wire v$FLOAT_4604_out0;
wire v$FLOAT_7676_out0;
wire v$FLOAT_7677_out0;
wire v$G10_10694_out0;
wire v$G10_10711_out0;
wire v$G10_130_out0;
wire v$G10_131_out0;
wire v$G10_13215_out0;
wire v$G10_13216_out0;
wire v$G10_13217_out0;
wire v$G10_13218_out0;
wire v$G10_1755_out0;
wire v$G10_1756_out0;
wire v$G10_1943_out0;
wire v$G10_1944_out0;
wire v$G10_1945_out0;
wire v$G10_1946_out0;
wire v$G10_2632_out0;
wire v$G10_2633_out0;
wire v$G10_2640_out0;
wire v$G10_2641_out0;
wire v$G10_2642_out0;
wire v$G10_2643_out0;
wire v$G10_4479_out0;
wire v$G10_4480_out0;
wire v$G10_602_out0;
wire v$G10_6975_out0;
wire v$G10_6976_out0;
wire v$G10_6977_out0;
wire v$G10_6978_out0;
wire v$G10_6979_out0;
wire v$G10_6980_out0;
wire v$G10_6981_out0;
wire v$G10_6982_out0;
wire v$G10_6983_out0;
wire v$G10_6984_out0;
wire v$G10_6985_out0;
wire v$G10_6986_out0;
wire v$G10_6987_out0;
wire v$G10_6988_out0;
wire v$G10_6989_out0;
wire v$G10_6990_out0;
wire v$G10_6991_out0;
wire v$G10_6992_out0;
wire v$G10_6993_out0;
wire v$G10_6994_out0;
wire v$G10_6995_out0;
wire v$G10_6996_out0;
wire v$G10_6997_out0;
wire v$G10_6998_out0;
wire v$G10_6999_out0;
wire v$G10_7000_out0;
wire v$G10_7001_out0;
wire v$G10_7002_out0;
wire v$G10_7003_out0;
wire v$G10_7004_out0;
wire v$G11_11165_out0;
wire v$G11_11166_out0;
wire v$G11_13342_out0;
wire v$G11_13343_out0;
wire v$G11_13344_out0;
wire v$G11_13345_out0;
wire v$G11_13439_out0;
wire v$G11_13440_out0;
wire v$G11_2550_out0;
wire v$G11_2551_out0;
wire v$G11_2626_out0;
wire v$G11_2627_out0;
wire v$G11_2937_out0;
wire v$G11_2938_out0;
wire v$G11_2939_out0;
wire v$G11_2940_out0;
wire v$G11_651_out0;
wire v$G11_652_out0;
wire v$G11_653_out0;
wire v$G11_654_out0;
wire v$G11_655_out0;
wire v$G11_656_out0;
wire v$G11_657_out0;
wire v$G11_658_out0;
wire v$G11_659_out0;
wire v$G11_660_out0;
wire v$G11_661_out0;
wire v$G11_662_out0;
wire v$G11_663_out0;
wire v$G11_664_out0;
wire v$G11_665_out0;
wire v$G11_666_out0;
wire v$G11_667_out0;
wire v$G11_668_out0;
wire v$G11_669_out0;
wire v$G11_670_out0;
wire v$G11_671_out0;
wire v$G11_672_out0;
wire v$G11_673_out0;
wire v$G11_674_out0;
wire v$G11_675_out0;
wire v$G11_676_out0;
wire v$G11_677_out0;
wire v$G11_678_out0;
wire v$G11_679_out0;
wire v$G11_680_out0;
wire v$G11_8652_out0;
wire v$G12_10321_out0;
wire v$G12_10322_out0;
wire v$G12_10688_out0;
wire v$G12_10689_out0;
wire v$G12_10690_out0;
wire v$G12_10691_out0;
wire v$G12_13221_out0;
wire v$G12_13222_out0;
wire v$G12_13223_out0;
wire v$G12_13224_out0;
wire v$G12_13225_out0;
wire v$G12_13226_out0;
wire v$G12_13227_out0;
wire v$G12_13228_out0;
wire v$G12_13229_out0;
wire v$G12_13230_out0;
wire v$G12_13231_out0;
wire v$G12_13232_out0;
wire v$G12_13233_out0;
wire v$G12_13234_out0;
wire v$G12_13235_out0;
wire v$G12_13236_out0;
wire v$G12_13237_out0;
wire v$G12_13238_out0;
wire v$G12_13239_out0;
wire v$G12_13240_out0;
wire v$G12_13241_out0;
wire v$G12_13242_out0;
wire v$G12_13243_out0;
wire v$G12_13244_out0;
wire v$G12_13245_out0;
wire v$G12_13246_out0;
wire v$G12_13247_out0;
wire v$G12_13248_out0;
wire v$G12_13249_out0;
wire v$G12_13250_out0;
wire v$G12_2270_out0;
wire v$G12_3345_out0;
wire v$G12_3346_out0;
wire v$G12_3347_out0;
wire v$G12_3348_out0;
wire v$G12_4699_out0;
wire v$G12_4700_out0;
wire v$G13_13352_out0;
wire v$G13_13353_out0;
wire v$G13_13354_out0;
wire v$G13_13355_out0;
wire v$G13_13356_out0;
wire v$G13_13357_out0;
wire v$G13_13358_out0;
wire v$G13_13359_out0;
wire v$G13_13360_out0;
wire v$G13_13361_out0;
wire v$G13_13362_out0;
wire v$G13_13363_out0;
wire v$G13_13364_out0;
wire v$G13_13365_out0;
wire v$G13_13366_out0;
wire v$G13_13367_out0;
wire v$G13_13368_out0;
wire v$G13_13369_out0;
wire v$G13_13370_out0;
wire v$G13_13371_out0;
wire v$G13_13372_out0;
wire v$G13_13373_out0;
wire v$G13_13374_out0;
wire v$G13_13375_out0;
wire v$G13_13376_out0;
wire v$G13_13377_out0;
wire v$G13_13378_out0;
wire v$G13_13379_out0;
wire v$G13_13380_out0;
wire v$G13_13381_out0;
wire v$G13_4705_out0;
wire v$G13_4706_out0;
wire v$G13_4707_out0;
wire v$G13_4708_out0;
wire v$G13_642_out0;
wire v$G13_643_out0;
wire v$G13_644_out0;
wire v$G13_645_out0;
wire v$G13_7083_out0;
wire v$G13_7084_out0;
wire v$G14_10407_out0;
wire v$G14_10408_out0;
wire v$G14_1178_out0;
wire v$G14_1179_out0;
wire v$G14_13268_out0;
wire v$G14_13269_out0;
wire v$G14_13672_out0;
wire v$G14_13673_out0;
wire v$G14_13674_out0;
wire v$G14_13675_out0;
wire v$G14_13676_out0;
wire v$G14_13677_out0;
wire v$G14_13678_out0;
wire v$G14_13679_out0;
wire v$G14_13680_out0;
wire v$G14_13681_out0;
wire v$G14_13682_out0;
wire v$G14_13683_out0;
wire v$G14_13684_out0;
wire v$G14_13685_out0;
wire v$G14_13686_out0;
wire v$G14_13687_out0;
wire v$G14_13688_out0;
wire v$G14_13689_out0;
wire v$G14_13690_out0;
wire v$G14_13691_out0;
wire v$G14_13692_out0;
wire v$G14_13693_out0;
wire v$G14_13694_out0;
wire v$G14_13695_out0;
wire v$G14_13696_out0;
wire v$G14_13697_out0;
wire v$G14_13698_out0;
wire v$G14_13699_out0;
wire v$G14_13700_out0;
wire v$G14_13701_out0;
wire v$G14_4533_out0;
wire v$G14_4534_out0;
wire v$G14_4535_out0;
wire v$G14_4536_out0;
wire v$G14_615_out0;
wire v$G14_616_out0;
wire v$G14_617_out0;
wire v$G14_618_out0;
wire v$G15_132_out0;
wire v$G15_133_out0;
wire v$G15_134_out0;
wire v$G15_135_out0;
wire v$G15_136_out0;
wire v$G15_137_out0;
wire v$G15_138_out0;
wire v$G15_139_out0;
wire v$G15_140_out0;
wire v$G15_141_out0;
wire v$G15_142_out0;
wire v$G15_143_out0;
wire v$G15_144_out0;
wire v$G15_145_out0;
wire v$G15_146_out0;
wire v$G15_147_out0;
wire v$G15_148_out0;
wire v$G15_149_out0;
wire v$G15_150_out0;
wire v$G15_151_out0;
wire v$G15_152_out0;
wire v$G15_153_out0;
wire v$G15_154_out0;
wire v$G15_155_out0;
wire v$G15_156_out0;
wire v$G15_157_out0;
wire v$G15_158_out0;
wire v$G15_159_out0;
wire v$G15_160_out0;
wire v$G15_161_out0;
wire v$G15_1814_out0;
wire v$G15_1815_out0;
wire v$G15_1816_out0;
wire v$G15_1817_out0;
wire v$G15_1855_out0;
wire v$G15_1856_out0;
wire v$G15_4654_out0;
wire v$G15_4655_out0;
wire v$G15_4656_out0;
wire v$G15_4657_out0;
wire v$G16_10906_out0;
wire v$G16_10907_out0;
wire v$G16_10908_out0;
wire v$G16_10909_out0;
wire v$G16_11034_out0;
wire v$G16_11035_out0;
wire v$G16_11036_out0;
wire v$G16_11037_out0;
wire v$G16_13183_out0;
wire v$G16_13184_out0;
wire v$G16_13185_out0;
wire v$G16_13186_out0;
wire v$G16_13187_out0;
wire v$G16_13188_out0;
wire v$G16_13189_out0;
wire v$G16_13190_out0;
wire v$G16_13191_out0;
wire v$G16_13192_out0;
wire v$G16_13193_out0;
wire v$G16_13194_out0;
wire v$G16_13195_out0;
wire v$G16_13196_out0;
wire v$G16_13197_out0;
wire v$G16_13198_out0;
wire v$G16_13199_out0;
wire v$G16_13200_out0;
wire v$G16_13201_out0;
wire v$G16_13202_out0;
wire v$G16_13203_out0;
wire v$G16_13204_out0;
wire v$G16_13205_out0;
wire v$G16_13206_out0;
wire v$G16_13207_out0;
wire v$G16_13208_out0;
wire v$G16_13209_out0;
wire v$G16_13210_out0;
wire v$G16_13211_out0;
wire v$G16_13212_out0;
wire v$G16_13388_out0;
wire v$G16_13389_out0;
wire v$G16_2310_out0;
wire v$G16_2311_out0;
wire v$G16_3024_out0;
wire v$G16_7701_out0;
wire v$G17_10710_out0;
wire v$G17_1903_out0;
wire v$G18_10489_out0;
wire v$G18_11204_out0;
wire v$G18_11205_out0;
wire v$G18_2407_out0;
wire v$G18_2408_out0;
wire v$G18_567_out0;
wire v$G18_8799_out0;
wire v$G18_8800_out0;
wire v$G18_8801_out0;
wire v$G18_8802_out0;
wire v$G19_10327_out0;
wire v$G19_10328_out0;
wire v$G19_3860_out0;
wire v$G19_4663_out0;
wire v$G19_4664_out0;
wire v$G1_10476_out0;
wire v$G1_10477_out0;
wire v$G1_10478_out0;
wire v$G1_10757_out0;
wire v$G1_10758_out0;
wire v$G1_10810_out0;
wire v$G1_11157_out0;
wire v$G1_11158_out0;
wire v$G1_1167_out0;
wire v$G1_1168_out0;
wire v$G1_1191_out0;
wire v$G1_1192_out0;
wire v$G1_13757_out0;
wire v$G1_13758_out0;
wire v$G1_13759_out0;
wire v$G1_13760_out0;
wire v$G1_13776_out0;
wire v$G1_13777_out0;
wire v$G1_1879_out0;
wire v$G1_1880_out0;
wire v$G1_1881_out0;
wire v$G1_1882_out0;
wire v$G1_1909_out0;
wire v$G1_1910_out0;
wire v$G1_1911_out0;
wire v$G1_1912_out0;
wire v$G1_1913_out0;
wire v$G1_1914_out0;
wire v$G1_1915_out0;
wire v$G1_1916_out0;
wire v$G1_1917_out0;
wire v$G1_1918_out0;
wire v$G1_1919_out0;
wire v$G1_1920_out0;
wire v$G1_1921_out0;
wire v$G1_1922_out0;
wire v$G1_1923_out0;
wire v$G1_1924_out0;
wire v$G1_1925_out0;
wire v$G1_1926_out0;
wire v$G1_1927_out0;
wire v$G1_1928_out0;
wire v$G1_1929_out0;
wire v$G1_1930_out0;
wire v$G1_1931_out0;
wire v$G1_1932_out0;
wire v$G1_1933_out0;
wire v$G1_1934_out0;
wire v$G1_1935_out0;
wire v$G1_1936_out0;
wire v$G1_1937_out0;
wire v$G1_1938_out0;
wire v$G1_2225_out0;
wire v$G1_2226_out0;
wire v$G1_2354_out0;
wire v$G1_2700_out0;
wire v$G1_2701_out0;
wire v$G1_2702_out0;
wire v$G1_2703_out0;
wire v$G1_2704_out0;
wire v$G1_2705_out0;
wire v$G1_2706_out0;
wire v$G1_2707_out0;
wire v$G1_2708_out0;
wire v$G1_2709_out0;
wire v$G1_2710_out0;
wire v$G1_2711_out0;
wire v$G1_2712_out0;
wire v$G1_2713_out0;
wire v$G1_2714_out0;
wire v$G1_2715_out0;
wire v$G1_277_out0;
wire v$G1_289_out0;
wire v$G1_290_out0;
wire v$G1_2911_out0;
wire v$G1_3018_out0;
wire v$G1_3019_out0;
wire v$G1_3995_out0;
wire v$G1_3996_out0;
wire v$G1_3997_out0;
wire v$G1_3998_out0;
wire v$G1_3999_out0;
wire v$G1_4000_out0;
wire v$G1_4001_out0;
wire v$G1_4002_out0;
wire v$G1_4003_out0;
wire v$G1_4004_out0;
wire v$G1_4005_out0;
wire v$G1_4006_out0;
wire v$G1_4007_out0;
wire v$G1_4008_out0;
wire v$G1_4009_out0;
wire v$G1_4010_out0;
wire v$G1_4011_out0;
wire v$G1_4012_out0;
wire v$G1_4013_out0;
wire v$G1_4014_out0;
wire v$G1_4015_out0;
wire v$G1_4016_out0;
wire v$G1_4017_out0;
wire v$G1_4018_out0;
wire v$G1_4019_out0;
wire v$G1_4020_out0;
wire v$G1_4021_out0;
wire v$G1_4022_out0;
wire v$G1_4023_out0;
wire v$G1_4024_out0;
wire v$G1_4025_out0;
wire v$G1_4026_out0;
wire v$G1_4027_out0;
wire v$G1_4028_out0;
wire v$G1_4029_out0;
wire v$G1_4030_out0;
wire v$G1_4031_out0;
wire v$G1_4032_out0;
wire v$G1_4033_out0;
wire v$G1_4034_out0;
wire v$G1_4035_out0;
wire v$G1_4036_out0;
wire v$G1_4037_out0;
wire v$G1_4038_out0;
wire v$G1_4039_out0;
wire v$G1_4040_out0;
wire v$G1_4041_out0;
wire v$G1_4042_out0;
wire v$G1_4043_out0;
wire v$G1_4044_out0;
wire v$G1_4045_out0;
wire v$G1_4046_out0;
wire v$G1_4047_out0;
wire v$G1_4048_out0;
wire v$G1_4049_out0;
wire v$G1_4050_out0;
wire v$G1_4051_out0;
wire v$G1_4052_out0;
wire v$G1_4053_out0;
wire v$G1_4054_out0;
wire v$G1_4055_out0;
wire v$G1_4056_out0;
wire v$G1_4057_out0;
wire v$G1_4058_out0;
wire v$G1_4059_out0;
wire v$G1_4060_out0;
wire v$G1_4061_out0;
wire v$G1_4062_out0;
wire v$G1_4063_out0;
wire v$G1_4064_out0;
wire v$G1_4065_out0;
wire v$G1_4066_out0;
wire v$G1_4067_out0;
wire v$G1_4068_out0;
wire v$G1_4069_out0;
wire v$G1_4070_out0;
wire v$G1_4071_out0;
wire v$G1_4072_out0;
wire v$G1_4073_out0;
wire v$G1_4074_out0;
wire v$G1_4075_out0;
wire v$G1_4076_out0;
wire v$G1_4077_out0;
wire v$G1_4078_out0;
wire v$G1_4079_out0;
wire v$G1_4080_out0;
wire v$G1_4081_out0;
wire v$G1_4082_out0;
wire v$G1_4083_out0;
wire v$G1_4084_out0;
wire v$G1_4085_out0;
wire v$G1_4086_out0;
wire v$G1_4087_out0;
wire v$G1_4088_out0;
wire v$G1_4089_out0;
wire v$G1_4090_out0;
wire v$G1_4091_out0;
wire v$G1_4092_out0;
wire v$G1_4093_out0;
wire v$G1_4094_out0;
wire v$G1_4095_out0;
wire v$G1_4096_out0;
wire v$G1_4097_out0;
wire v$G1_4098_out0;
wire v$G1_4099_out0;
wire v$G1_4100_out0;
wire v$G1_4101_out0;
wire v$G1_4102_out0;
wire v$G1_4103_out0;
wire v$G1_4104_out0;
wire v$G1_4105_out0;
wire v$G1_4106_out0;
wire v$G1_4107_out0;
wire v$G1_4108_out0;
wire v$G1_4109_out0;
wire v$G1_4110_out0;
wire v$G1_4111_out0;
wire v$G1_4112_out0;
wire v$G1_4113_out0;
wire v$G1_4114_out0;
wire v$G1_4115_out0;
wire v$G1_4116_out0;
wire v$G1_4117_out0;
wire v$G1_4118_out0;
wire v$G1_4119_out0;
wire v$G1_4120_out0;
wire v$G1_4121_out0;
wire v$G1_4122_out0;
wire v$G1_4123_out0;
wire v$G1_4124_out0;
wire v$G1_4125_out0;
wire v$G1_4126_out0;
wire v$G1_4127_out0;
wire v$G1_4128_out0;
wire v$G1_4129_out0;
wire v$G1_4130_out0;
wire v$G1_4131_out0;
wire v$G1_4132_out0;
wire v$G1_4133_out0;
wire v$G1_4134_out0;
wire v$G1_4135_out0;
wire v$G1_4136_out0;
wire v$G1_4137_out0;
wire v$G1_4138_out0;
wire v$G1_4139_out0;
wire v$G1_4140_out0;
wire v$G1_4141_out0;
wire v$G1_4142_out0;
wire v$G1_4143_out0;
wire v$G1_4144_out0;
wire v$G1_4145_out0;
wire v$G1_4146_out0;
wire v$G1_4147_out0;
wire v$G1_4148_out0;
wire v$G1_4149_out0;
wire v$G1_4150_out0;
wire v$G1_4151_out0;
wire v$G1_4152_out0;
wire v$G1_4153_out0;
wire v$G1_4154_out0;
wire v$G1_4155_out0;
wire v$G1_4156_out0;
wire v$G1_4157_out0;
wire v$G1_4158_out0;
wire v$G1_4159_out0;
wire v$G1_4160_out0;
wire v$G1_4161_out0;
wire v$G1_4162_out0;
wire v$G1_4163_out0;
wire v$G1_4164_out0;
wire v$G1_4165_out0;
wire v$G1_4166_out0;
wire v$G1_4167_out0;
wire v$G1_4168_out0;
wire v$G1_4169_out0;
wire v$G1_4170_out0;
wire v$G1_4171_out0;
wire v$G1_4172_out0;
wire v$G1_4173_out0;
wire v$G1_4174_out0;
wire v$G1_4175_out0;
wire v$G1_4176_out0;
wire v$G1_4177_out0;
wire v$G1_4178_out0;
wire v$G1_4179_out0;
wire v$G1_4180_out0;
wire v$G1_4181_out0;
wire v$G1_4182_out0;
wire v$G1_4183_out0;
wire v$G1_4184_out0;
wire v$G1_4185_out0;
wire v$G1_4186_out0;
wire v$G1_4187_out0;
wire v$G1_4188_out0;
wire v$G1_4189_out0;
wire v$G1_4190_out0;
wire v$G1_4191_out0;
wire v$G1_4192_out0;
wire v$G1_4193_out0;
wire v$G1_4194_out0;
wire v$G1_4195_out0;
wire v$G1_4196_out0;
wire v$G1_4197_out0;
wire v$G1_4198_out0;
wire v$G1_4199_out0;
wire v$G1_4200_out0;
wire v$G1_4201_out0;
wire v$G1_4202_out0;
wire v$G1_4203_out0;
wire v$G1_4204_out0;
wire v$G1_4205_out0;
wire v$G1_4206_out0;
wire v$G1_4207_out0;
wire v$G1_4208_out0;
wire v$G1_4209_out0;
wire v$G1_4210_out0;
wire v$G1_4211_out0;
wire v$G1_4212_out0;
wire v$G1_4213_out0;
wire v$G1_4214_out0;
wire v$G1_4215_out0;
wire v$G1_4216_out0;
wire v$G1_4217_out0;
wire v$G1_4218_out0;
wire v$G1_4219_out0;
wire v$G1_4220_out0;
wire v$G1_4221_out0;
wire v$G1_4222_out0;
wire v$G1_4223_out0;
wire v$G1_4224_out0;
wire v$G1_4225_out0;
wire v$G1_4226_out0;
wire v$G1_4227_out0;
wire v$G1_4228_out0;
wire v$G1_4229_out0;
wire v$G1_4230_out0;
wire v$G1_4231_out0;
wire v$G1_4232_out0;
wire v$G1_4233_out0;
wire v$G1_4234_out0;
wire v$G1_4235_out0;
wire v$G1_4236_out0;
wire v$G1_4237_out0;
wire v$G1_4238_out0;
wire v$G1_4239_out0;
wire v$G1_4240_out0;
wire v$G1_4241_out0;
wire v$G1_4242_out0;
wire v$G1_4243_out0;
wire v$G1_4244_out0;
wire v$G1_4245_out0;
wire v$G1_4246_out0;
wire v$G1_4247_out0;
wire v$G1_4248_out0;
wire v$G1_4249_out0;
wire v$G1_4250_out0;
wire v$G1_4251_out0;
wire v$G1_4252_out0;
wire v$G1_4253_out0;
wire v$G1_4254_out0;
wire v$G1_4255_out0;
wire v$G1_4256_out0;
wire v$G1_4257_out0;
wire v$G1_4258_out0;
wire v$G1_4259_out0;
wire v$G1_4260_out0;
wire v$G1_4261_out0;
wire v$G1_4262_out0;
wire v$G1_4263_out0;
wire v$G1_4264_out0;
wire v$G1_4265_out0;
wire v$G1_4266_out0;
wire v$G1_4267_out0;
wire v$G1_4268_out0;
wire v$G1_4269_out0;
wire v$G1_4270_out0;
wire v$G1_4271_out0;
wire v$G1_4272_out0;
wire v$G1_4273_out0;
wire v$G1_4274_out0;
wire v$G1_4275_out0;
wire v$G1_4276_out0;
wire v$G1_4277_out0;
wire v$G1_4278_out0;
wire v$G1_4279_out0;
wire v$G1_4280_out0;
wire v$G1_4281_out0;
wire v$G1_4282_out0;
wire v$G1_4283_out0;
wire v$G1_4284_out0;
wire v$G1_4285_out0;
wire v$G1_4286_out0;
wire v$G1_4287_out0;
wire v$G1_4288_out0;
wire v$G1_4289_out0;
wire v$G1_4290_out0;
wire v$G1_4291_out0;
wire v$G1_4292_out0;
wire v$G1_4293_out0;
wire v$G1_4294_out0;
wire v$G1_4295_out0;
wire v$G1_4296_out0;
wire v$G1_4297_out0;
wire v$G1_4298_out0;
wire v$G1_4299_out0;
wire v$G1_4300_out0;
wire v$G1_4301_out0;
wire v$G1_4302_out0;
wire v$G1_4303_out0;
wire v$G1_4304_out0;
wire v$G1_4305_out0;
wire v$G1_4306_out0;
wire v$G1_4307_out0;
wire v$G1_4308_out0;
wire v$G1_4309_out0;
wire v$G1_4310_out0;
wire v$G1_4311_out0;
wire v$G1_4312_out0;
wire v$G1_4313_out0;
wire v$G1_4314_out0;
wire v$G1_4315_out0;
wire v$G1_4316_out0;
wire v$G1_4317_out0;
wire v$G1_4318_out0;
wire v$G1_4319_out0;
wire v$G1_4320_out0;
wire v$G1_4321_out0;
wire v$G1_4322_out0;
wire v$G1_4323_out0;
wire v$G1_4324_out0;
wire v$G1_4325_out0;
wire v$G1_4326_out0;
wire v$G1_4327_out0;
wire v$G1_4328_out0;
wire v$G1_4329_out0;
wire v$G1_4330_out0;
wire v$G1_4331_out0;
wire v$G1_4332_out0;
wire v$G1_4333_out0;
wire v$G1_4334_out0;
wire v$G1_4335_out0;
wire v$G1_4336_out0;
wire v$G1_4337_out0;
wire v$G1_4338_out0;
wire v$G1_4339_out0;
wire v$G1_4340_out0;
wire v$G1_4341_out0;
wire v$G1_4342_out0;
wire v$G1_4343_out0;
wire v$G1_4344_out0;
wire v$G1_4345_out0;
wire v$G1_4346_out0;
wire v$G1_4347_out0;
wire v$G1_4348_out0;
wire v$G1_4349_out0;
wire v$G1_4350_out0;
wire v$G1_4351_out0;
wire v$G1_4352_out0;
wire v$G1_4353_out0;
wire v$G1_4354_out0;
wire v$G1_4355_out0;
wire v$G1_4356_out0;
wire v$G1_4357_out0;
wire v$G1_4358_out0;
wire v$G1_4359_out0;
wire v$G1_4360_out0;
wire v$G1_4361_out0;
wire v$G1_4362_out0;
wire v$G1_4363_out0;
wire v$G1_4364_out0;
wire v$G1_4365_out0;
wire v$G1_4366_out0;
wire v$G1_4367_out0;
wire v$G1_4368_out0;
wire v$G1_4369_out0;
wire v$G1_4370_out0;
wire v$G1_4371_out0;
wire v$G1_4372_out0;
wire v$G1_4373_out0;
wire v$G1_4374_out0;
wire v$G1_4375_out0;
wire v$G1_4376_out0;
wire v$G1_4377_out0;
wire v$G1_4378_out0;
wire v$G1_4379_out0;
wire v$G1_4380_out0;
wire v$G1_4381_out0;
wire v$G1_4382_out0;
wire v$G1_4383_out0;
wire v$G1_4384_out0;
wire v$G1_4385_out0;
wire v$G1_4386_out0;
wire v$G1_4387_out0;
wire v$G1_4388_out0;
wire v$G1_4389_out0;
wire v$G1_4390_out0;
wire v$G1_4391_out0;
wire v$G1_4392_out0;
wire v$G1_4393_out0;
wire v$G1_4394_out0;
wire v$G1_4395_out0;
wire v$G1_4396_out0;
wire v$G1_4397_out0;
wire v$G1_4398_out0;
wire v$G1_4399_out0;
wire v$G1_4400_out0;
wire v$G1_4401_out0;
wire v$G1_4402_out0;
wire v$G1_4403_out0;
wire v$G1_4404_out0;
wire v$G1_4405_out0;
wire v$G1_4406_out0;
wire v$G1_4407_out0;
wire v$G1_4408_out0;
wire v$G1_4409_out0;
wire v$G1_4410_out0;
wire v$G1_4411_out0;
wire v$G1_4412_out0;
wire v$G1_4413_out0;
wire v$G1_4414_out0;
wire v$G1_4415_out0;
wire v$G1_4416_out0;
wire v$G1_4417_out0;
wire v$G1_4418_out0;
wire v$G1_4419_out0;
wire v$G1_4420_out0;
wire v$G1_4421_out0;
wire v$G1_4422_out0;
wire v$G1_4423_out0;
wire v$G1_4424_out0;
wire v$G1_4425_out0;
wire v$G1_4426_out0;
wire v$G1_4427_out0;
wire v$G1_4428_out0;
wire v$G1_4429_out0;
wire v$G1_4430_out0;
wire v$G1_4431_out0;
wire v$G1_4432_out0;
wire v$G1_4433_out0;
wire v$G1_4434_out0;
wire v$G1_4435_out0;
wire v$G1_4436_out0;
wire v$G1_4437_out0;
wire v$G1_4438_out0;
wire v$G1_4439_out0;
wire v$G1_4440_out0;
wire v$G1_4441_out0;
wire v$G1_4442_out0;
wire v$G1_646_out0;
wire v$G1_647_out0;
wire v$G1_7717_out0;
wire v$G1_7718_out0;
wire v$G1_7719_out0;
wire v$G1_7720_out0;
wire v$G1_7721_out0;
wire v$G1_7722_out0;
wire v$G1_7723_out0;
wire v$G1_7724_out0;
wire v$G1_7725_out0;
wire v$G1_7726_out0;
wire v$G1_7727_out0;
wire v$G1_7728_out0;
wire v$G1_7729_out0;
wire v$G1_7730_out0;
wire v$G1_7731_out0;
wire v$G1_7732_out0;
wire v$G1_7733_out0;
wire v$G1_7734_out0;
wire v$G1_7735_out0;
wire v$G1_7736_out0;
wire v$G1_7737_out0;
wire v$G1_7738_out0;
wire v$G1_7739_out0;
wire v$G1_7740_out0;
wire v$G1_7741_out0;
wire v$G1_7742_out0;
wire v$G1_7743_out0;
wire v$G1_7744_out0;
wire v$G1_7745_out0;
wire v$G1_7746_out0;
wire v$G1_7747_out0;
wire v$G1_7748_out0;
wire v$G1_7749_out0;
wire v$G1_7750_out0;
wire v$G1_7751_out0;
wire v$G1_7752_out0;
wire v$G1_7753_out0;
wire v$G1_7754_out0;
wire v$G1_7755_out0;
wire v$G1_7756_out0;
wire v$G1_7757_out0;
wire v$G1_7758_out0;
wire v$G1_7759_out0;
wire v$G1_7760_out0;
wire v$G1_7761_out0;
wire v$G1_7762_out0;
wire v$G1_7763_out0;
wire v$G1_7764_out0;
wire v$G1_7765_out0;
wire v$G1_7766_out0;
wire v$G1_7767_out0;
wire v$G1_7768_out0;
wire v$G1_7769_out0;
wire v$G1_7770_out0;
wire v$G1_7771_out0;
wire v$G1_7772_out0;
wire v$G1_7773_out0;
wire v$G1_7774_out0;
wire v$G1_7775_out0;
wire v$G1_7776_out0;
wire v$G1_7777_out0;
wire v$G1_7778_out0;
wire v$G1_7779_out0;
wire v$G1_7780_out0;
wire v$G1_7781_out0;
wire v$G1_7782_out0;
wire v$G1_7783_out0;
wire v$G1_7784_out0;
wire v$G1_7785_out0;
wire v$G1_7786_out0;
wire v$G1_7787_out0;
wire v$G1_7788_out0;
wire v$G1_7789_out0;
wire v$G1_7790_out0;
wire v$G1_7791_out0;
wire v$G1_7792_out0;
wire v$G1_7793_out0;
wire v$G1_7794_out0;
wire v$G1_7795_out0;
wire v$G1_7796_out0;
wire v$G1_7797_out0;
wire v$G1_7798_out0;
wire v$G1_7799_out0;
wire v$G1_7800_out0;
wire v$G1_7801_out0;
wire v$G1_7802_out0;
wire v$G1_7803_out0;
wire v$G1_7804_out0;
wire v$G1_7805_out0;
wire v$G1_7806_out0;
wire v$G1_7807_out0;
wire v$G1_7808_out0;
wire v$G1_7809_out0;
wire v$G1_7810_out0;
wire v$G1_7811_out0;
wire v$G1_7812_out0;
wire v$G1_7813_out0;
wire v$G1_7814_out0;
wire v$G1_7815_out0;
wire v$G1_7816_out0;
wire v$G1_7817_out0;
wire v$G1_7818_out0;
wire v$G1_7819_out0;
wire v$G1_7820_out0;
wire v$G1_7821_out0;
wire v$G1_7822_out0;
wire v$G1_7823_out0;
wire v$G1_7824_out0;
wire v$G1_7825_out0;
wire v$G1_7826_out0;
wire v$G1_7827_out0;
wire v$G1_7828_out0;
wire v$G1_7829_out0;
wire v$G1_7830_out0;
wire v$G1_7831_out0;
wire v$G1_7832_out0;
wire v$G1_7833_out0;
wire v$G1_7834_out0;
wire v$G1_7835_out0;
wire v$G1_7836_out0;
wire v$G1_7837_out0;
wire v$G1_7838_out0;
wire v$G1_7839_out0;
wire v$G1_7840_out0;
wire v$G1_7841_out0;
wire v$G1_7842_out0;
wire v$G1_7843_out0;
wire v$G1_7844_out0;
wire v$G1_7845_out0;
wire v$G1_7846_out0;
wire v$G1_7847_out0;
wire v$G1_7848_out0;
wire v$G1_7849_out0;
wire v$G1_7850_out0;
wire v$G1_7851_out0;
wire v$G1_7852_out0;
wire v$G1_7853_out0;
wire v$G1_7854_out0;
wire v$G1_7855_out0;
wire v$G1_7856_out0;
wire v$G1_7857_out0;
wire v$G1_7858_out0;
wire v$G1_7859_out0;
wire v$G1_7860_out0;
wire v$G1_7861_out0;
wire v$G1_7862_out0;
wire v$G1_7863_out0;
wire v$G1_7864_out0;
wire v$G1_7865_out0;
wire v$G1_7866_out0;
wire v$G1_7867_out0;
wire v$G1_7868_out0;
wire v$G1_7869_out0;
wire v$G1_7870_out0;
wire v$G1_7871_out0;
wire v$G1_7872_out0;
wire v$G1_7873_out0;
wire v$G1_7874_out0;
wire v$G1_7875_out0;
wire v$G1_7876_out0;
wire v$G1_7877_out0;
wire v$G1_7878_out0;
wire v$G1_7879_out0;
wire v$G1_7880_out0;
wire v$G1_7881_out0;
wire v$G1_7882_out0;
wire v$G1_7883_out0;
wire v$G1_7884_out0;
wire v$G1_7885_out0;
wire v$G1_7886_out0;
wire v$G1_7887_out0;
wire v$G1_7888_out0;
wire v$G1_7889_out0;
wire v$G1_7890_out0;
wire v$G1_7891_out0;
wire v$G1_7892_out0;
wire v$G1_7893_out0;
wire v$G1_7894_out0;
wire v$G1_7895_out0;
wire v$G1_7896_out0;
wire v$G1_7897_out0;
wire v$G1_7898_out0;
wire v$G1_7899_out0;
wire v$G1_7900_out0;
wire v$G1_7901_out0;
wire v$G1_7902_out0;
wire v$G1_7903_out0;
wire v$G1_7904_out0;
wire v$G1_7905_out0;
wire v$G1_7906_out0;
wire v$G1_7907_out0;
wire v$G1_7908_out0;
wire v$G1_7909_out0;
wire v$G1_7910_out0;
wire v$G1_7911_out0;
wire v$G1_7912_out0;
wire v$G1_7913_out0;
wire v$G1_7914_out0;
wire v$G1_7915_out0;
wire v$G1_7916_out0;
wire v$G1_7917_out0;
wire v$G1_7918_out0;
wire v$G1_7919_out0;
wire v$G1_7920_out0;
wire v$G1_7921_out0;
wire v$G1_7922_out0;
wire v$G1_7923_out0;
wire v$G1_7924_out0;
wire v$G1_7925_out0;
wire v$G1_7926_out0;
wire v$G1_7927_out0;
wire v$G1_7928_out0;
wire v$G1_7929_out0;
wire v$G1_7930_out0;
wire v$G1_7931_out0;
wire v$G1_7932_out0;
wire v$G1_7933_out0;
wire v$G1_7934_out0;
wire v$G1_7935_out0;
wire v$G1_7936_out0;
wire v$G1_7937_out0;
wire v$G1_7938_out0;
wire v$G1_7939_out0;
wire v$G1_7940_out0;
wire v$G1_7941_out0;
wire v$G1_7942_out0;
wire v$G1_7943_out0;
wire v$G1_7944_out0;
wire v$G1_7945_out0;
wire v$G1_7946_out0;
wire v$G1_7947_out0;
wire v$G1_7948_out0;
wire v$G1_7949_out0;
wire v$G1_7950_out0;
wire v$G1_7951_out0;
wire v$G1_7952_out0;
wire v$G1_7953_out0;
wire v$G1_7954_out0;
wire v$G1_7955_out0;
wire v$G1_7956_out0;
wire v$G1_7957_out0;
wire v$G1_7958_out0;
wire v$G1_7959_out0;
wire v$G1_7960_out0;
wire v$G1_7961_out0;
wire v$G1_7962_out0;
wire v$G1_7963_out0;
wire v$G1_7964_out0;
wire v$G1_7965_out0;
wire v$G1_7966_out0;
wire v$G1_7967_out0;
wire v$G1_7968_out0;
wire v$G1_7969_out0;
wire v$G1_7970_out0;
wire v$G1_7971_out0;
wire v$G1_7972_out0;
wire v$G1_7973_out0;
wire v$G1_7974_out0;
wire v$G1_7975_out0;
wire v$G1_7976_out0;
wire v$G1_7977_out0;
wire v$G1_7978_out0;
wire v$G1_7979_out0;
wire v$G1_7980_out0;
wire v$G1_7981_out0;
wire v$G1_7982_out0;
wire v$G1_7983_out0;
wire v$G1_7984_out0;
wire v$G1_7985_out0;
wire v$G1_7986_out0;
wire v$G1_7987_out0;
wire v$G1_7988_out0;
wire v$G1_7989_out0;
wire v$G1_7990_out0;
wire v$G1_7991_out0;
wire v$G1_7992_out0;
wire v$G1_7993_out0;
wire v$G1_7994_out0;
wire v$G1_7995_out0;
wire v$G1_7996_out0;
wire v$G1_7997_out0;
wire v$G1_7998_out0;
wire v$G1_7999_out0;
wire v$G1_8000_out0;
wire v$G1_8001_out0;
wire v$G1_8002_out0;
wire v$G1_8003_out0;
wire v$G1_8004_out0;
wire v$G1_8005_out0;
wire v$G1_8006_out0;
wire v$G1_8007_out0;
wire v$G1_8008_out0;
wire v$G1_8009_out0;
wire v$G1_8010_out0;
wire v$G1_8011_out0;
wire v$G1_8012_out0;
wire v$G1_8013_out0;
wire v$G1_8014_out0;
wire v$G1_8015_out0;
wire v$G1_8016_out0;
wire v$G1_8017_out0;
wire v$G1_8018_out0;
wire v$G1_8019_out0;
wire v$G1_8020_out0;
wire v$G1_8021_out0;
wire v$G1_8022_out0;
wire v$G1_8023_out0;
wire v$G1_8024_out0;
wire v$G1_8025_out0;
wire v$G1_8026_out0;
wire v$G1_8027_out0;
wire v$G1_8028_out0;
wire v$G1_8029_out0;
wire v$G1_8030_out0;
wire v$G1_8031_out0;
wire v$G1_8032_out0;
wire v$G1_8033_out0;
wire v$G1_8034_out0;
wire v$G1_8035_out0;
wire v$G1_8036_out0;
wire v$G1_8037_out0;
wire v$G1_8038_out0;
wire v$G1_8039_out0;
wire v$G1_8040_out0;
wire v$G1_8041_out0;
wire v$G1_8042_out0;
wire v$G1_8043_out0;
wire v$G1_8044_out0;
wire v$G1_8045_out0;
wire v$G1_8046_out0;
wire v$G1_8047_out0;
wire v$G1_8048_out0;
wire v$G1_8049_out0;
wire v$G1_8050_out0;
wire v$G1_8051_out0;
wire v$G1_8052_out0;
wire v$G1_8053_out0;
wire v$G1_8054_out0;
wire v$G1_8055_out0;
wire v$G1_8056_out0;
wire v$G1_8057_out0;
wire v$G1_8058_out0;
wire v$G1_8059_out0;
wire v$G1_8060_out0;
wire v$G1_8061_out0;
wire v$G1_8062_out0;
wire v$G1_8063_out0;
wire v$G1_8064_out0;
wire v$G1_8065_out0;
wire v$G1_8066_out0;
wire v$G1_8067_out0;
wire v$G1_8068_out0;
wire v$G1_8069_out0;
wire v$G1_8070_out0;
wire v$G1_8071_out0;
wire v$G1_8072_out0;
wire v$G1_8073_out0;
wire v$G1_8074_out0;
wire v$G1_8075_out0;
wire v$G1_8076_out0;
wire v$G1_8077_out0;
wire v$G1_8078_out0;
wire v$G1_8079_out0;
wire v$G1_8080_out0;
wire v$G1_8081_out0;
wire v$G1_8082_out0;
wire v$G1_8083_out0;
wire v$G1_8084_out0;
wire v$G1_8085_out0;
wire v$G1_8086_out0;
wire v$G1_8087_out0;
wire v$G1_8088_out0;
wire v$G1_8089_out0;
wire v$G1_8090_out0;
wire v$G1_8091_out0;
wire v$G1_8092_out0;
wire v$G1_8093_out0;
wire v$G1_8094_out0;
wire v$G1_8095_out0;
wire v$G1_8096_out0;
wire v$G1_8097_out0;
wire v$G1_8098_out0;
wire v$G1_8099_out0;
wire v$G1_8100_out0;
wire v$G1_8101_out0;
wire v$G1_8102_out0;
wire v$G1_8103_out0;
wire v$G1_8104_out0;
wire v$G1_8105_out0;
wire v$G1_8106_out0;
wire v$G1_8107_out0;
wire v$G1_8108_out0;
wire v$G1_8109_out0;
wire v$G1_8110_out0;
wire v$G1_8111_out0;
wire v$G1_8112_out0;
wire v$G1_8113_out0;
wire v$G1_8114_out0;
wire v$G1_8115_out0;
wire v$G1_8116_out0;
wire v$G1_8117_out0;
wire v$G1_8118_out0;
wire v$G1_8119_out0;
wire v$G1_8120_out0;
wire v$G1_8121_out0;
wire v$G1_8122_out0;
wire v$G1_8123_out0;
wire v$G1_8124_out0;
wire v$G1_8125_out0;
wire v$G1_8126_out0;
wire v$G1_8127_out0;
wire v$G1_8128_out0;
wire v$G1_8129_out0;
wire v$G1_8130_out0;
wire v$G1_8131_out0;
wire v$G1_8132_out0;
wire v$G1_8133_out0;
wire v$G1_8134_out0;
wire v$G1_8135_out0;
wire v$G1_8136_out0;
wire v$G1_8137_out0;
wire v$G1_8138_out0;
wire v$G1_8139_out0;
wire v$G1_8140_out0;
wire v$G1_8141_out0;
wire v$G1_8142_out0;
wire v$G1_8143_out0;
wire v$G1_8144_out0;
wire v$G1_8145_out0;
wire v$G1_8146_out0;
wire v$G1_8147_out0;
wire v$G1_8148_out0;
wire v$G1_8149_out0;
wire v$G1_8150_out0;
wire v$G1_8151_out0;
wire v$G1_8152_out0;
wire v$G1_8153_out0;
wire v$G1_8154_out0;
wire v$G1_8155_out0;
wire v$G1_8156_out0;
wire v$G1_8157_out0;
wire v$G1_8158_out0;
wire v$G1_8159_out0;
wire v$G1_8160_out0;
wire v$G1_8161_out0;
wire v$G1_8162_out0;
wire v$G1_8163_out0;
wire v$G1_8164_out0;
wire v$G1_8165_out0;
wire v$G1_8166_out0;
wire v$G1_8167_out0;
wire v$G1_8168_out0;
wire v$G1_8169_out0;
wire v$G1_8170_out0;
wire v$G1_8171_out0;
wire v$G1_8172_out0;
wire v$G1_8173_out0;
wire v$G1_8174_out0;
wire v$G1_8175_out0;
wire v$G1_8176_out0;
wire v$G1_8177_out0;
wire v$G1_8178_out0;
wire v$G1_8179_out0;
wire v$G1_8180_out0;
wire v$G1_8181_out0;
wire v$G1_8182_out0;
wire v$G1_8183_out0;
wire v$G1_8184_out0;
wire v$G1_8185_out0;
wire v$G1_8186_out0;
wire v$G1_8187_out0;
wire v$G1_8188_out0;
wire v$G1_8189_out0;
wire v$G1_8190_out0;
wire v$G1_8191_out0;
wire v$G1_8192_out0;
wire v$G1_8193_out0;
wire v$G1_8194_out0;
wire v$G1_8195_out0;
wire v$G1_8196_out0;
wire v$G1_8197_out0;
wire v$G1_8198_out0;
wire v$G1_8199_out0;
wire v$G1_8200_out0;
wire v$G1_8201_out0;
wire v$G1_8202_out0;
wire v$G1_8203_out0;
wire v$G1_8204_out0;
wire v$G1_8205_out0;
wire v$G1_8206_out0;
wire v$G1_8207_out0;
wire v$G1_8208_out0;
wire v$G1_8209_out0;
wire v$G1_8210_out0;
wire v$G1_8211_out0;
wire v$G1_8212_out0;
wire v$G1_8213_out0;
wire v$G1_8214_out0;
wire v$G1_8215_out0;
wire v$G1_8216_out0;
wire v$G1_8217_out0;
wire v$G1_8218_out0;
wire v$G1_8219_out0;
wire v$G1_8220_out0;
wire v$G1_8221_out0;
wire v$G1_8222_out0;
wire v$G1_8223_out0;
wire v$G1_8224_out0;
wire v$G1_8225_out0;
wire v$G1_8226_out0;
wire v$G1_8227_out0;
wire v$G1_8228_out0;
wire v$G1_8229_out0;
wire v$G1_8230_out0;
wire v$G1_8231_out0;
wire v$G1_8232_out0;
wire v$G1_8233_out0;
wire v$G1_8234_out0;
wire v$G1_8235_out0;
wire v$G1_8236_out0;
wire v$G1_8237_out0;
wire v$G1_8238_out0;
wire v$G1_8239_out0;
wire v$G1_8240_out0;
wire v$G1_8241_out0;
wire v$G1_8242_out0;
wire v$G1_8243_out0;
wire v$G1_8244_out0;
wire v$G1_8245_out0;
wire v$G1_8246_out0;
wire v$G1_8247_out0;
wire v$G1_8248_out0;
wire v$G1_8249_out0;
wire v$G1_8250_out0;
wire v$G1_8251_out0;
wire v$G1_8252_out0;
wire v$G1_8253_out0;
wire v$G1_8254_out0;
wire v$G1_8255_out0;
wire v$G1_8256_out0;
wire v$G1_8257_out0;
wire v$G1_8258_out0;
wire v$G1_8259_out0;
wire v$G1_8260_out0;
wire v$G1_8261_out0;
wire v$G1_8262_out0;
wire v$G1_8263_out0;
wire v$G1_8264_out0;
wire v$G1_8265_out0;
wire v$G1_8266_out0;
wire v$G1_8267_out0;
wire v$G1_8268_out0;
wire v$G1_8269_out0;
wire v$G1_8270_out0;
wire v$G1_8271_out0;
wire v$G1_8272_out0;
wire v$G1_8273_out0;
wire v$G1_8274_out0;
wire v$G1_8275_out0;
wire v$G1_8276_out0;
wire v$G1_8277_out0;
wire v$G1_8278_out0;
wire v$G1_8279_out0;
wire v$G1_8280_out0;
wire v$G1_8281_out0;
wire v$G1_8282_out0;
wire v$G1_8283_out0;
wire v$G1_8284_out0;
wire v$G1_8285_out0;
wire v$G1_8286_out0;
wire v$G1_8287_out0;
wire v$G1_8288_out0;
wire v$G1_8289_out0;
wire v$G1_8290_out0;
wire v$G1_8291_out0;
wire v$G1_8292_out0;
wire v$G1_8293_out0;
wire v$G1_8294_out0;
wire v$G1_8295_out0;
wire v$G1_8296_out0;
wire v$G1_8297_out0;
wire v$G1_8298_out0;
wire v$G1_8299_out0;
wire v$G1_8300_out0;
wire v$G1_8301_out0;
wire v$G1_8302_out0;
wire v$G1_8303_out0;
wire v$G1_8304_out0;
wire v$G1_8305_out0;
wire v$G1_8306_out0;
wire v$G1_8307_out0;
wire v$G1_8308_out0;
wire v$G1_8309_out0;
wire v$G1_8310_out0;
wire v$G1_8311_out0;
wire v$G1_8312_out0;
wire v$G1_8313_out0;
wire v$G1_8314_out0;
wire v$G1_8315_out0;
wire v$G1_8316_out0;
wire v$G1_8317_out0;
wire v$G1_8318_out0;
wire v$G1_8319_out0;
wire v$G1_8320_out0;
wire v$G1_8321_out0;
wire v$G1_8322_out0;
wire v$G1_8323_out0;
wire v$G1_8324_out0;
wire v$G1_8325_out0;
wire v$G1_8326_out0;
wire v$G1_8327_out0;
wire v$G1_8328_out0;
wire v$G1_8329_out0;
wire v$G1_8330_out0;
wire v$G1_8331_out0;
wire v$G1_8332_out0;
wire v$G1_8333_out0;
wire v$G1_8334_out0;
wire v$G1_8335_out0;
wire v$G1_8336_out0;
wire v$G1_8337_out0;
wire v$G1_8338_out0;
wire v$G1_8339_out0;
wire v$G1_8340_out0;
wire v$G1_8341_out0;
wire v$G1_8342_out0;
wire v$G1_8343_out0;
wire v$G1_8344_out0;
wire v$G1_8345_out0;
wire v$G1_8346_out0;
wire v$G1_8347_out0;
wire v$G1_8348_out0;
wire v$G1_8349_out0;
wire v$G1_8350_out0;
wire v$G1_8351_out0;
wire v$G1_8352_out0;
wire v$G1_8353_out0;
wire v$G1_8354_out0;
wire v$G1_8355_out0;
wire v$G1_8356_out0;
wire v$G1_8357_out0;
wire v$G1_8358_out0;
wire v$G1_8359_out0;
wire v$G1_8360_out0;
wire v$G1_8361_out0;
wire v$G1_8362_out0;
wire v$G1_8363_out0;
wire v$G1_8364_out0;
wire v$G1_8365_out0;
wire v$G1_8366_out0;
wire v$G1_8367_out0;
wire v$G1_8368_out0;
wire v$G1_8369_out0;
wire v$G1_8370_out0;
wire v$G1_8371_out0;
wire v$G1_8372_out0;
wire v$G1_8373_out0;
wire v$G1_8374_out0;
wire v$G1_8375_out0;
wire v$G1_8376_out0;
wire v$G1_8377_out0;
wire v$G1_8378_out0;
wire v$G1_8379_out0;
wire v$G1_8380_out0;
wire v$G1_8381_out0;
wire v$G1_8382_out0;
wire v$G1_8383_out0;
wire v$G1_8384_out0;
wire v$G1_8385_out0;
wire v$G1_8386_out0;
wire v$G1_8387_out0;
wire v$G1_8388_out0;
wire v$G1_8389_out0;
wire v$G1_8390_out0;
wire v$G1_8391_out0;
wire v$G1_8392_out0;
wire v$G1_8393_out0;
wire v$G1_8394_out0;
wire v$G1_8395_out0;
wire v$G1_8396_out0;
wire v$G1_8397_out0;
wire v$G1_8398_out0;
wire v$G1_8399_out0;
wire v$G1_8400_out0;
wire v$G1_8401_out0;
wire v$G1_8402_out0;
wire v$G1_8403_out0;
wire v$G1_8404_out0;
wire v$G1_8405_out0;
wire v$G1_8406_out0;
wire v$G1_8407_out0;
wire v$G1_8408_out0;
wire v$G1_8409_out0;
wire v$G1_8410_out0;
wire v$G1_8411_out0;
wire v$G1_8412_out0;
wire v$G1_8413_out0;
wire v$G1_8414_out0;
wire v$G1_8415_out0;
wire v$G1_8416_out0;
wire v$G1_8417_out0;
wire v$G1_8418_out0;
wire v$G1_8419_out0;
wire v$G1_8420_out0;
wire v$G1_8421_out0;
wire v$G1_8422_out0;
wire v$G1_8423_out0;
wire v$G1_8424_out0;
wire v$G1_8425_out0;
wire v$G1_8426_out0;
wire v$G1_8427_out0;
wire v$G1_8428_out0;
wire v$G1_8429_out0;
wire v$G1_8430_out0;
wire v$G1_8431_out0;
wire v$G1_8432_out0;
wire v$G1_8433_out0;
wire v$G1_8434_out0;
wire v$G1_8435_out0;
wire v$G1_8436_out0;
wire v$G1_8437_out0;
wire v$G1_8438_out0;
wire v$G1_8439_out0;
wire v$G1_8440_out0;
wire v$G1_8441_out0;
wire v$G1_8442_out0;
wire v$G1_8443_out0;
wire v$G1_8444_out0;
wire v$G1_8445_out0;
wire v$G1_8446_out0;
wire v$G1_8447_out0;
wire v$G1_8448_out0;
wire v$G1_8449_out0;
wire v$G1_8450_out0;
wire v$G1_8451_out0;
wire v$G1_8452_out0;
wire v$G1_8453_out0;
wire v$G1_8454_out0;
wire v$G1_8455_out0;
wire v$G1_8456_out0;
wire v$G1_8457_out0;
wire v$G1_8458_out0;
wire v$G1_8459_out0;
wire v$G1_8460_out0;
wire v$G1_8461_out0;
wire v$G1_8462_out0;
wire v$G1_8463_out0;
wire v$G1_8464_out0;
wire v$G1_8465_out0;
wire v$G1_8466_out0;
wire v$G1_8467_out0;
wire v$G1_8468_out0;
wire v$G1_8469_out0;
wire v$G1_8470_out0;
wire v$G1_8471_out0;
wire v$G1_8472_out0;
wire v$G1_8473_out0;
wire v$G1_8474_out0;
wire v$G1_8475_out0;
wire v$G1_8476_out0;
wire v$G1_8477_out0;
wire v$G1_8478_out0;
wire v$G1_8479_out0;
wire v$G1_8480_out0;
wire v$G1_8481_out0;
wire v$G1_8482_out0;
wire v$G1_8483_out0;
wire v$G1_8484_out0;
wire v$G1_8485_out0;
wire v$G1_8486_out0;
wire v$G1_8487_out0;
wire v$G1_8488_out0;
wire v$G1_8489_out0;
wire v$G1_8490_out0;
wire v$G1_8491_out0;
wire v$G1_8492_out0;
wire v$G1_8493_out0;
wire v$G1_8494_out0;
wire v$G1_8495_out0;
wire v$G1_8496_out0;
wire v$G1_8497_out0;
wire v$G1_8498_out0;
wire v$G1_8499_out0;
wire v$G1_8500_out0;
wire v$G1_8501_out0;
wire v$G1_8502_out0;
wire v$G1_8503_out0;
wire v$G1_8504_out0;
wire v$G1_8505_out0;
wire v$G1_8506_out0;
wire v$G1_8507_out0;
wire v$G1_8508_out0;
wire v$G1_8509_out0;
wire v$G1_8510_out0;
wire v$G1_8511_out0;
wire v$G1_8512_out0;
wire v$G1_8513_out0;
wire v$G1_8514_out0;
wire v$G1_8515_out0;
wire v$G1_8516_out0;
wire v$G1_8517_out0;
wire v$G1_8518_out0;
wire v$G1_8519_out0;
wire v$G1_8520_out0;
wire v$G1_8521_out0;
wire v$G1_8522_out0;
wire v$G1_8523_out0;
wire v$G1_8524_out0;
wire v$G1_8525_out0;
wire v$G1_8526_out0;
wire v$G1_8527_out0;
wire v$G1_8528_out0;
wire v$G1_8529_out0;
wire v$G1_8530_out0;
wire v$G1_8531_out0;
wire v$G1_8532_out0;
wire v$G1_8533_out0;
wire v$G1_8534_out0;
wire v$G1_8535_out0;
wire v$G1_8536_out0;
wire v$G1_8537_out0;
wire v$G1_8538_out0;
wire v$G1_8539_out0;
wire v$G1_8540_out0;
wire v$G1_8541_out0;
wire v$G1_8542_out0;
wire v$G1_8543_out0;
wire v$G1_8544_out0;
wire v$G1_8545_out0;
wire v$G1_8546_out0;
wire v$G1_8547_out0;
wire v$G1_8548_out0;
wire v$G1_8549_out0;
wire v$G1_8550_out0;
wire v$G1_8551_out0;
wire v$G1_8552_out0;
wire v$G1_8553_out0;
wire v$G1_8554_out0;
wire v$G1_8555_out0;
wire v$G1_8556_out0;
wire v$G1_8557_out0;
wire v$G1_8558_out0;
wire v$G1_8559_out0;
wire v$G1_8560_out0;
wire v$G1_8561_out0;
wire v$G1_8562_out0;
wire v$G1_8563_out0;
wire v$G1_8564_out0;
wire v$G1_8565_out0;
wire v$G1_8566_out0;
wire v$G1_8567_out0;
wire v$G1_8568_out0;
wire v$G1_8569_out0;
wire v$G1_8570_out0;
wire v$G1_8571_out0;
wire v$G1_8572_out0;
wire v$G1_8573_out0;
wire v$G1_8574_out0;
wire v$G1_8575_out0;
wire v$G1_8576_out0;
wire v$G1_8577_out0;
wire v$G1_8578_out0;
wire v$G1_8579_out0;
wire v$G1_8580_out0;
wire v$G1_8581_out0;
wire v$G1_8582_out0;
wire v$G1_8583_out0;
wire v$G1_8584_out0;
wire v$G1_8585_out0;
wire v$G1_8586_out0;
wire v$G1_8587_out0;
wire v$G1_8588_out0;
wire v$G1_8589_out0;
wire v$G1_8590_out0;
wire v$G1_8591_out0;
wire v$G1_8592_out0;
wire v$G1_8593_out0;
wire v$G1_8594_out0;
wire v$G1_8595_out0;
wire v$G1_8596_out0;
wire v$G1_8597_out0;
wire v$G1_8598_out0;
wire v$G1_8599_out0;
wire v$G1_8600_out0;
wire v$G1_8601_out0;
wire v$G1_8602_out0;
wire v$G1_8603_out0;
wire v$G1_8604_out0;
wire v$G1_8605_out0;
wire v$G1_8606_out0;
wire v$G1_8607_out0;
wire v$G1_8608_out0;
wire v$G1_8609_out0;
wire v$G1_8610_out0;
wire v$G1_8611_out0;
wire v$G1_8612_out0;
wire v$G1_8613_out0;
wire v$G1_8614_out0;
wire v$G1_8615_out0;
wire v$G1_8616_out0;
wire v$G1_8617_out0;
wire v$G1_8618_out0;
wire v$G1_8619_out0;
wire v$G1_8620_out0;
wire v$G1_8621_out0;
wire v$G1_8622_out0;
wire v$G1_8623_out0;
wire v$G1_8624_out0;
wire v$G1_8625_out0;
wire v$G1_8626_out0;
wire v$G1_8627_out0;
wire v$G1_8628_out0;
wire v$G1_8629_out0;
wire v$G1_8630_out0;
wire v$G1_8631_out0;
wire v$G1_8632_out0;
wire v$G1_8633_out0;
wire v$G1_8634_out0;
wire v$G1_8635_out0;
wire v$G1_8636_out0;
wire v$G1_8637_out0;
wire v$G1_8638_out0;
wire v$G1_8639_out0;
wire v$G1_8640_out0;
wire v$G1_8641_out0;
wire v$G1_8642_out0;
wire v$G1_8643_out0;
wire v$G1_8644_out0;
wire v$G1_8693_out0;
wire v$G1_8694_out0;
wire v$G1_8695_out0;
wire v$G1_8696_out0;
wire v$G20_11040_out0;
wire v$G20_11147_out0;
wire v$G20_11148_out0;
wire v$G20_598_out0;
wire v$G20_599_out0;
wire v$G21_10681_out0;
wire v$G21_10788_out0;
wire v$G21_2656_out0;
wire v$G21_2657_out0;
wire v$G21_2885_out0;
wire v$G21_2886_out0;
wire v$G21_3808_out0;
wire v$G21_3809_out0;
wire v$G21_3810_out0;
wire v$G21_3811_out0;
wire v$G22_10620_out0;
wire v$G22_10983_out0;
wire v$G22_10984_out0;
wire v$G22_10985_out0;
wire v$G22_10986_out0;
wire v$G22_13663_out0;
wire v$G22_13707_out0;
wire v$G22_13708_out0;
wire v$G22_1899_out0;
wire v$G22_1900_out0;
wire v$G23_10439_out0;
wire v$G23_10440_out0;
wire v$G23_2614_out0;
wire v$G23_2840_out0;
wire v$G23_2841_out0;
wire v$G23_3083_out0;
wire v$G23_4852_out0;
wire v$G23_4853_out0;
wire v$G23_4854_out0;
wire v$G23_4855_out0;
wire v$G24_10460_out0;
wire v$G24_10560_out0;
wire v$G24_10561_out0;
wire v$G24_10562_out0;
wire v$G24_10563_out0;
wire v$G24_3955_out0;
wire v$G24_3956_out0;
wire v$G24_4780_out0;
wire v$G25_4658_out0;
wire v$G25_6962_out0;
wire v$G25_6963_out0;
wire v$G26_4735_out0;
wire v$G26_4736_out0;
wire v$G27_9793_out0;
wire v$G27_9794_out0;
wire v$G28_2098_out0;
wire v$G28_2099_out0;
wire v$G28_2100_out0;
wire v$G28_2101_out0;
wire v$G28_6868_out0;
wire v$G28_6869_out0;
wire v$G29_5834_out0;
wire v$G29_5835_out0;
wire v$G2_10278_out0;
wire v$G2_10471_out0;
wire v$G2_10799_out0;
wire v$G2_10800_out0;
wire v$G2_11134_out0;
wire v$G2_11135_out0;
wire v$G2_12230_out0;
wire v$G2_12231_out0;
wire v$G2_12253_out0;
wire v$G2_12254_out0;
wire v$G2_12255_out0;
wire v$G2_12256_out0;
wire v$G2_12257_out0;
wire v$G2_12258_out0;
wire v$G2_12259_out0;
wire v$G2_12260_out0;
wire v$G2_12261_out0;
wire v$G2_12262_out0;
wire v$G2_12263_out0;
wire v$G2_12264_out0;
wire v$G2_12265_out0;
wire v$G2_12266_out0;
wire v$G2_12267_out0;
wire v$G2_12268_out0;
wire v$G2_12269_out0;
wire v$G2_12270_out0;
wire v$G2_12271_out0;
wire v$G2_12272_out0;
wire v$G2_12273_out0;
wire v$G2_12274_out0;
wire v$G2_12275_out0;
wire v$G2_12276_out0;
wire v$G2_12277_out0;
wire v$G2_12278_out0;
wire v$G2_12279_out0;
wire v$G2_12280_out0;
wire v$G2_12281_out0;
wire v$G2_12282_out0;
wire v$G2_12283_out0;
wire v$G2_12284_out0;
wire v$G2_12285_out0;
wire v$G2_12286_out0;
wire v$G2_12287_out0;
wire v$G2_12288_out0;
wire v$G2_12289_out0;
wire v$G2_12290_out0;
wire v$G2_12291_out0;
wire v$G2_12292_out0;
wire v$G2_12293_out0;
wire v$G2_12294_out0;
wire v$G2_12295_out0;
wire v$G2_12296_out0;
wire v$G2_12297_out0;
wire v$G2_12298_out0;
wire v$G2_12299_out0;
wire v$G2_12300_out0;
wire v$G2_12301_out0;
wire v$G2_12302_out0;
wire v$G2_12303_out0;
wire v$G2_12304_out0;
wire v$G2_12305_out0;
wire v$G2_12306_out0;
wire v$G2_12307_out0;
wire v$G2_12308_out0;
wire v$G2_12309_out0;
wire v$G2_12310_out0;
wire v$G2_12311_out0;
wire v$G2_12312_out0;
wire v$G2_12313_out0;
wire v$G2_12314_out0;
wire v$G2_12315_out0;
wire v$G2_12316_out0;
wire v$G2_12317_out0;
wire v$G2_12318_out0;
wire v$G2_12319_out0;
wire v$G2_12320_out0;
wire v$G2_12321_out0;
wire v$G2_12322_out0;
wire v$G2_12323_out0;
wire v$G2_12324_out0;
wire v$G2_12325_out0;
wire v$G2_12326_out0;
wire v$G2_12327_out0;
wire v$G2_12328_out0;
wire v$G2_12329_out0;
wire v$G2_12330_out0;
wire v$G2_12331_out0;
wire v$G2_12332_out0;
wire v$G2_12333_out0;
wire v$G2_12334_out0;
wire v$G2_12335_out0;
wire v$G2_12336_out0;
wire v$G2_12337_out0;
wire v$G2_12338_out0;
wire v$G2_12339_out0;
wire v$G2_12340_out0;
wire v$G2_12341_out0;
wire v$G2_12342_out0;
wire v$G2_12343_out0;
wire v$G2_12344_out0;
wire v$G2_12345_out0;
wire v$G2_12346_out0;
wire v$G2_12347_out0;
wire v$G2_12348_out0;
wire v$G2_12349_out0;
wire v$G2_12350_out0;
wire v$G2_12351_out0;
wire v$G2_12352_out0;
wire v$G2_12353_out0;
wire v$G2_12354_out0;
wire v$G2_12355_out0;
wire v$G2_12356_out0;
wire v$G2_12357_out0;
wire v$G2_12358_out0;
wire v$G2_12359_out0;
wire v$G2_12360_out0;
wire v$G2_12361_out0;
wire v$G2_12362_out0;
wire v$G2_12363_out0;
wire v$G2_12364_out0;
wire v$G2_12365_out0;
wire v$G2_12366_out0;
wire v$G2_12367_out0;
wire v$G2_12368_out0;
wire v$G2_12369_out0;
wire v$G2_12370_out0;
wire v$G2_12371_out0;
wire v$G2_12372_out0;
wire v$G2_12373_out0;
wire v$G2_12374_out0;
wire v$G2_12375_out0;
wire v$G2_12376_out0;
wire v$G2_12377_out0;
wire v$G2_12378_out0;
wire v$G2_12379_out0;
wire v$G2_12380_out0;
wire v$G2_12381_out0;
wire v$G2_12382_out0;
wire v$G2_12383_out0;
wire v$G2_12384_out0;
wire v$G2_12385_out0;
wire v$G2_12386_out0;
wire v$G2_12387_out0;
wire v$G2_12388_out0;
wire v$G2_12389_out0;
wire v$G2_12390_out0;
wire v$G2_12391_out0;
wire v$G2_12392_out0;
wire v$G2_12393_out0;
wire v$G2_12394_out0;
wire v$G2_12395_out0;
wire v$G2_12396_out0;
wire v$G2_12397_out0;
wire v$G2_12398_out0;
wire v$G2_12399_out0;
wire v$G2_12400_out0;
wire v$G2_12401_out0;
wire v$G2_12402_out0;
wire v$G2_12403_out0;
wire v$G2_12404_out0;
wire v$G2_12405_out0;
wire v$G2_12406_out0;
wire v$G2_12407_out0;
wire v$G2_12408_out0;
wire v$G2_12409_out0;
wire v$G2_12410_out0;
wire v$G2_12411_out0;
wire v$G2_12412_out0;
wire v$G2_12413_out0;
wire v$G2_12414_out0;
wire v$G2_12415_out0;
wire v$G2_12416_out0;
wire v$G2_12417_out0;
wire v$G2_12418_out0;
wire v$G2_12419_out0;
wire v$G2_12420_out0;
wire v$G2_12421_out0;
wire v$G2_12422_out0;
wire v$G2_12423_out0;
wire v$G2_12424_out0;
wire v$G2_12425_out0;
wire v$G2_12426_out0;
wire v$G2_12427_out0;
wire v$G2_12428_out0;
wire v$G2_12429_out0;
wire v$G2_12430_out0;
wire v$G2_12431_out0;
wire v$G2_12432_out0;
wire v$G2_12433_out0;
wire v$G2_12434_out0;
wire v$G2_12435_out0;
wire v$G2_12436_out0;
wire v$G2_12437_out0;
wire v$G2_12438_out0;
wire v$G2_12439_out0;
wire v$G2_12440_out0;
wire v$G2_12441_out0;
wire v$G2_12442_out0;
wire v$G2_12443_out0;
wire v$G2_12444_out0;
wire v$G2_12445_out0;
wire v$G2_12446_out0;
wire v$G2_12447_out0;
wire v$G2_12448_out0;
wire v$G2_12449_out0;
wire v$G2_12450_out0;
wire v$G2_12451_out0;
wire v$G2_12452_out0;
wire v$G2_12453_out0;
wire v$G2_12454_out0;
wire v$G2_12455_out0;
wire v$G2_12456_out0;
wire v$G2_12457_out0;
wire v$G2_12458_out0;
wire v$G2_12459_out0;
wire v$G2_12460_out0;
wire v$G2_12461_out0;
wire v$G2_12462_out0;
wire v$G2_12463_out0;
wire v$G2_12464_out0;
wire v$G2_12465_out0;
wire v$G2_12466_out0;
wire v$G2_12467_out0;
wire v$G2_12468_out0;
wire v$G2_12469_out0;
wire v$G2_12470_out0;
wire v$G2_12471_out0;
wire v$G2_12472_out0;
wire v$G2_12473_out0;
wire v$G2_12474_out0;
wire v$G2_12475_out0;
wire v$G2_12476_out0;
wire v$G2_12477_out0;
wire v$G2_12478_out0;
wire v$G2_12479_out0;
wire v$G2_12480_out0;
wire v$G2_12481_out0;
wire v$G2_12482_out0;
wire v$G2_12483_out0;
wire v$G2_12484_out0;
wire v$G2_12485_out0;
wire v$G2_12486_out0;
wire v$G2_12487_out0;
wire v$G2_12488_out0;
wire v$G2_12489_out0;
wire v$G2_12490_out0;
wire v$G2_12491_out0;
wire v$G2_12492_out0;
wire v$G2_12493_out0;
wire v$G2_12494_out0;
wire v$G2_12495_out0;
wire v$G2_12496_out0;
wire v$G2_12497_out0;
wire v$G2_12498_out0;
wire v$G2_12499_out0;
wire v$G2_12500_out0;
wire v$G2_12501_out0;
wire v$G2_12502_out0;
wire v$G2_12503_out0;
wire v$G2_12504_out0;
wire v$G2_12505_out0;
wire v$G2_12506_out0;
wire v$G2_12507_out0;
wire v$G2_12508_out0;
wire v$G2_12509_out0;
wire v$G2_12510_out0;
wire v$G2_12511_out0;
wire v$G2_12512_out0;
wire v$G2_12513_out0;
wire v$G2_12514_out0;
wire v$G2_12515_out0;
wire v$G2_12516_out0;
wire v$G2_12517_out0;
wire v$G2_12518_out0;
wire v$G2_12519_out0;
wire v$G2_12520_out0;
wire v$G2_12521_out0;
wire v$G2_12522_out0;
wire v$G2_12523_out0;
wire v$G2_12524_out0;
wire v$G2_12525_out0;
wire v$G2_12526_out0;
wire v$G2_12527_out0;
wire v$G2_12528_out0;
wire v$G2_12529_out0;
wire v$G2_12530_out0;
wire v$G2_12531_out0;
wire v$G2_12532_out0;
wire v$G2_12533_out0;
wire v$G2_12534_out0;
wire v$G2_12535_out0;
wire v$G2_12536_out0;
wire v$G2_12537_out0;
wire v$G2_12538_out0;
wire v$G2_12539_out0;
wire v$G2_12540_out0;
wire v$G2_12541_out0;
wire v$G2_12542_out0;
wire v$G2_12543_out0;
wire v$G2_12544_out0;
wire v$G2_12545_out0;
wire v$G2_12546_out0;
wire v$G2_12547_out0;
wire v$G2_12548_out0;
wire v$G2_12549_out0;
wire v$G2_12550_out0;
wire v$G2_12551_out0;
wire v$G2_12552_out0;
wire v$G2_12553_out0;
wire v$G2_12554_out0;
wire v$G2_12555_out0;
wire v$G2_12556_out0;
wire v$G2_12557_out0;
wire v$G2_12558_out0;
wire v$G2_12559_out0;
wire v$G2_12560_out0;
wire v$G2_12561_out0;
wire v$G2_12562_out0;
wire v$G2_12563_out0;
wire v$G2_12564_out0;
wire v$G2_12565_out0;
wire v$G2_12566_out0;
wire v$G2_12567_out0;
wire v$G2_12568_out0;
wire v$G2_12569_out0;
wire v$G2_12570_out0;
wire v$G2_12571_out0;
wire v$G2_12572_out0;
wire v$G2_12573_out0;
wire v$G2_12574_out0;
wire v$G2_12575_out0;
wire v$G2_12576_out0;
wire v$G2_12577_out0;
wire v$G2_12578_out0;
wire v$G2_12579_out0;
wire v$G2_12580_out0;
wire v$G2_12581_out0;
wire v$G2_12582_out0;
wire v$G2_12583_out0;
wire v$G2_12584_out0;
wire v$G2_12585_out0;
wire v$G2_12586_out0;
wire v$G2_12587_out0;
wire v$G2_12588_out0;
wire v$G2_12589_out0;
wire v$G2_12590_out0;
wire v$G2_12591_out0;
wire v$G2_12592_out0;
wire v$G2_12593_out0;
wire v$G2_12594_out0;
wire v$G2_12595_out0;
wire v$G2_12596_out0;
wire v$G2_12597_out0;
wire v$G2_12598_out0;
wire v$G2_12599_out0;
wire v$G2_12600_out0;
wire v$G2_12601_out0;
wire v$G2_12602_out0;
wire v$G2_12603_out0;
wire v$G2_12604_out0;
wire v$G2_12605_out0;
wire v$G2_12606_out0;
wire v$G2_12607_out0;
wire v$G2_12608_out0;
wire v$G2_12609_out0;
wire v$G2_12610_out0;
wire v$G2_12611_out0;
wire v$G2_12612_out0;
wire v$G2_12613_out0;
wire v$G2_12614_out0;
wire v$G2_12615_out0;
wire v$G2_12616_out0;
wire v$G2_12617_out0;
wire v$G2_12618_out0;
wire v$G2_12619_out0;
wire v$G2_12620_out0;
wire v$G2_12621_out0;
wire v$G2_12622_out0;
wire v$G2_12623_out0;
wire v$G2_12624_out0;
wire v$G2_12625_out0;
wire v$G2_12626_out0;
wire v$G2_12627_out0;
wire v$G2_12628_out0;
wire v$G2_12629_out0;
wire v$G2_12630_out0;
wire v$G2_12631_out0;
wire v$G2_12632_out0;
wire v$G2_12633_out0;
wire v$G2_12634_out0;
wire v$G2_12635_out0;
wire v$G2_12636_out0;
wire v$G2_12637_out0;
wire v$G2_12638_out0;
wire v$G2_12639_out0;
wire v$G2_12640_out0;
wire v$G2_12641_out0;
wire v$G2_12642_out0;
wire v$G2_12643_out0;
wire v$G2_12644_out0;
wire v$G2_12645_out0;
wire v$G2_12646_out0;
wire v$G2_12647_out0;
wire v$G2_12648_out0;
wire v$G2_12649_out0;
wire v$G2_12650_out0;
wire v$G2_12651_out0;
wire v$G2_12652_out0;
wire v$G2_12653_out0;
wire v$G2_12654_out0;
wire v$G2_12655_out0;
wire v$G2_12656_out0;
wire v$G2_12657_out0;
wire v$G2_12658_out0;
wire v$G2_12659_out0;
wire v$G2_12660_out0;
wire v$G2_12661_out0;
wire v$G2_12662_out0;
wire v$G2_12663_out0;
wire v$G2_12664_out0;
wire v$G2_12665_out0;
wire v$G2_12666_out0;
wire v$G2_12667_out0;
wire v$G2_12668_out0;
wire v$G2_12669_out0;
wire v$G2_12670_out0;
wire v$G2_12671_out0;
wire v$G2_12672_out0;
wire v$G2_12673_out0;
wire v$G2_12674_out0;
wire v$G2_12675_out0;
wire v$G2_12676_out0;
wire v$G2_12677_out0;
wire v$G2_12678_out0;
wire v$G2_12679_out0;
wire v$G2_12680_out0;
wire v$G2_12681_out0;
wire v$G2_12682_out0;
wire v$G2_12683_out0;
wire v$G2_12684_out0;
wire v$G2_12685_out0;
wire v$G2_12686_out0;
wire v$G2_12687_out0;
wire v$G2_12688_out0;
wire v$G2_12689_out0;
wire v$G2_12690_out0;
wire v$G2_12691_out0;
wire v$G2_12692_out0;
wire v$G2_12693_out0;
wire v$G2_12694_out0;
wire v$G2_12695_out0;
wire v$G2_12696_out0;
wire v$G2_12697_out0;
wire v$G2_12698_out0;
wire v$G2_12699_out0;
wire v$G2_12700_out0;
wire v$G2_12701_out0;
wire v$G2_12702_out0;
wire v$G2_12703_out0;
wire v$G2_12704_out0;
wire v$G2_12705_out0;
wire v$G2_12706_out0;
wire v$G2_12707_out0;
wire v$G2_12708_out0;
wire v$G2_12709_out0;
wire v$G2_12710_out0;
wire v$G2_12711_out0;
wire v$G2_12712_out0;
wire v$G2_12713_out0;
wire v$G2_12714_out0;
wire v$G2_12715_out0;
wire v$G2_12716_out0;
wire v$G2_12717_out0;
wire v$G2_12718_out0;
wire v$G2_12719_out0;
wire v$G2_12720_out0;
wire v$G2_12721_out0;
wire v$G2_12722_out0;
wire v$G2_12723_out0;
wire v$G2_12724_out0;
wire v$G2_12725_out0;
wire v$G2_12726_out0;
wire v$G2_12727_out0;
wire v$G2_12728_out0;
wire v$G2_12729_out0;
wire v$G2_12730_out0;
wire v$G2_12731_out0;
wire v$G2_12732_out0;
wire v$G2_12733_out0;
wire v$G2_12734_out0;
wire v$G2_12735_out0;
wire v$G2_12736_out0;
wire v$G2_12737_out0;
wire v$G2_12738_out0;
wire v$G2_12739_out0;
wire v$G2_12740_out0;
wire v$G2_12741_out0;
wire v$G2_12742_out0;
wire v$G2_12743_out0;
wire v$G2_12744_out0;
wire v$G2_12745_out0;
wire v$G2_12746_out0;
wire v$G2_12747_out0;
wire v$G2_12748_out0;
wire v$G2_12749_out0;
wire v$G2_12750_out0;
wire v$G2_12751_out0;
wire v$G2_12752_out0;
wire v$G2_12753_out0;
wire v$G2_12754_out0;
wire v$G2_12755_out0;
wire v$G2_12756_out0;
wire v$G2_12757_out0;
wire v$G2_12758_out0;
wire v$G2_12759_out0;
wire v$G2_12760_out0;
wire v$G2_12761_out0;
wire v$G2_12762_out0;
wire v$G2_12763_out0;
wire v$G2_12764_out0;
wire v$G2_12765_out0;
wire v$G2_12766_out0;
wire v$G2_12767_out0;
wire v$G2_12768_out0;
wire v$G2_12769_out0;
wire v$G2_12770_out0;
wire v$G2_12771_out0;
wire v$G2_12772_out0;
wire v$G2_12773_out0;
wire v$G2_12774_out0;
wire v$G2_12775_out0;
wire v$G2_12776_out0;
wire v$G2_12777_out0;
wire v$G2_12778_out0;
wire v$G2_12779_out0;
wire v$G2_12780_out0;
wire v$G2_12781_out0;
wire v$G2_12782_out0;
wire v$G2_12783_out0;
wire v$G2_12784_out0;
wire v$G2_12785_out0;
wire v$G2_12786_out0;
wire v$G2_12787_out0;
wire v$G2_12788_out0;
wire v$G2_12789_out0;
wire v$G2_12790_out0;
wire v$G2_12791_out0;
wire v$G2_12792_out0;
wire v$G2_12793_out0;
wire v$G2_12794_out0;
wire v$G2_12795_out0;
wire v$G2_12796_out0;
wire v$G2_12797_out0;
wire v$G2_12798_out0;
wire v$G2_12799_out0;
wire v$G2_12800_out0;
wire v$G2_12801_out0;
wire v$G2_12802_out0;
wire v$G2_12803_out0;
wire v$G2_12804_out0;
wire v$G2_12805_out0;
wire v$G2_12806_out0;
wire v$G2_12807_out0;
wire v$G2_12808_out0;
wire v$G2_12809_out0;
wire v$G2_12810_out0;
wire v$G2_12811_out0;
wire v$G2_12812_out0;
wire v$G2_12813_out0;
wire v$G2_12814_out0;
wire v$G2_12815_out0;
wire v$G2_12816_out0;
wire v$G2_12817_out0;
wire v$G2_12818_out0;
wire v$G2_12819_out0;
wire v$G2_12820_out0;
wire v$G2_12821_out0;
wire v$G2_12822_out0;
wire v$G2_12823_out0;
wire v$G2_12824_out0;
wire v$G2_12825_out0;
wire v$G2_12826_out0;
wire v$G2_12827_out0;
wire v$G2_12828_out0;
wire v$G2_12829_out0;
wire v$G2_12830_out0;
wire v$G2_12831_out0;
wire v$G2_12832_out0;
wire v$G2_12833_out0;
wire v$G2_12834_out0;
wire v$G2_12835_out0;
wire v$G2_12836_out0;
wire v$G2_12837_out0;
wire v$G2_12838_out0;
wire v$G2_12839_out0;
wire v$G2_12840_out0;
wire v$G2_12841_out0;
wire v$G2_12842_out0;
wire v$G2_12843_out0;
wire v$G2_12844_out0;
wire v$G2_12845_out0;
wire v$G2_12846_out0;
wire v$G2_12847_out0;
wire v$G2_12848_out0;
wire v$G2_12849_out0;
wire v$G2_12850_out0;
wire v$G2_12851_out0;
wire v$G2_12852_out0;
wire v$G2_12853_out0;
wire v$G2_12854_out0;
wire v$G2_12855_out0;
wire v$G2_12856_out0;
wire v$G2_12857_out0;
wire v$G2_12858_out0;
wire v$G2_12859_out0;
wire v$G2_12860_out0;
wire v$G2_12861_out0;
wire v$G2_12862_out0;
wire v$G2_12863_out0;
wire v$G2_12864_out0;
wire v$G2_12865_out0;
wire v$G2_12866_out0;
wire v$G2_12867_out0;
wire v$G2_12868_out0;
wire v$G2_12869_out0;
wire v$G2_12870_out0;
wire v$G2_12871_out0;
wire v$G2_12872_out0;
wire v$G2_12873_out0;
wire v$G2_12874_out0;
wire v$G2_12875_out0;
wire v$G2_12876_out0;
wire v$G2_12877_out0;
wire v$G2_12878_out0;
wire v$G2_12879_out0;
wire v$G2_12880_out0;
wire v$G2_12881_out0;
wire v$G2_12882_out0;
wire v$G2_12883_out0;
wire v$G2_12884_out0;
wire v$G2_12885_out0;
wire v$G2_12886_out0;
wire v$G2_12887_out0;
wire v$G2_12888_out0;
wire v$G2_12889_out0;
wire v$G2_12890_out0;
wire v$G2_12891_out0;
wire v$G2_12892_out0;
wire v$G2_12893_out0;
wire v$G2_12894_out0;
wire v$G2_12895_out0;
wire v$G2_12896_out0;
wire v$G2_12897_out0;
wire v$G2_12898_out0;
wire v$G2_12899_out0;
wire v$G2_12900_out0;
wire v$G2_12901_out0;
wire v$G2_12902_out0;
wire v$G2_12903_out0;
wire v$G2_12904_out0;
wire v$G2_12905_out0;
wire v$G2_12906_out0;
wire v$G2_12907_out0;
wire v$G2_12908_out0;
wire v$G2_12909_out0;
wire v$G2_12910_out0;
wire v$G2_12911_out0;
wire v$G2_12912_out0;
wire v$G2_12913_out0;
wire v$G2_12914_out0;
wire v$G2_12915_out0;
wire v$G2_12916_out0;
wire v$G2_12917_out0;
wire v$G2_12918_out0;
wire v$G2_12919_out0;
wire v$G2_12920_out0;
wire v$G2_12921_out0;
wire v$G2_12922_out0;
wire v$G2_12923_out0;
wire v$G2_12924_out0;
wire v$G2_12925_out0;
wire v$G2_12926_out0;
wire v$G2_12927_out0;
wire v$G2_12928_out0;
wire v$G2_12929_out0;
wire v$G2_12930_out0;
wire v$G2_12931_out0;
wire v$G2_12932_out0;
wire v$G2_12933_out0;
wire v$G2_12934_out0;
wire v$G2_12935_out0;
wire v$G2_12936_out0;
wire v$G2_12937_out0;
wire v$G2_12938_out0;
wire v$G2_12939_out0;
wire v$G2_12940_out0;
wire v$G2_12941_out0;
wire v$G2_12942_out0;
wire v$G2_12943_out0;
wire v$G2_12944_out0;
wire v$G2_12945_out0;
wire v$G2_12946_out0;
wire v$G2_12947_out0;
wire v$G2_12948_out0;
wire v$G2_12949_out0;
wire v$G2_12950_out0;
wire v$G2_12951_out0;
wire v$G2_12952_out0;
wire v$G2_12953_out0;
wire v$G2_12954_out0;
wire v$G2_12955_out0;
wire v$G2_12956_out0;
wire v$G2_12957_out0;
wire v$G2_12958_out0;
wire v$G2_12959_out0;
wire v$G2_12960_out0;
wire v$G2_12961_out0;
wire v$G2_12962_out0;
wire v$G2_12963_out0;
wire v$G2_12964_out0;
wire v$G2_12965_out0;
wire v$G2_12966_out0;
wire v$G2_12967_out0;
wire v$G2_12968_out0;
wire v$G2_12969_out0;
wire v$G2_12970_out0;
wire v$G2_12971_out0;
wire v$G2_12972_out0;
wire v$G2_12973_out0;
wire v$G2_12974_out0;
wire v$G2_12975_out0;
wire v$G2_12976_out0;
wire v$G2_12977_out0;
wire v$G2_12978_out0;
wire v$G2_12979_out0;
wire v$G2_12980_out0;
wire v$G2_12981_out0;
wire v$G2_12982_out0;
wire v$G2_12983_out0;
wire v$G2_12984_out0;
wire v$G2_12985_out0;
wire v$G2_12986_out0;
wire v$G2_12987_out0;
wire v$G2_12988_out0;
wire v$G2_12989_out0;
wire v$G2_12990_out0;
wire v$G2_12991_out0;
wire v$G2_12992_out0;
wire v$G2_12993_out0;
wire v$G2_12994_out0;
wire v$G2_12995_out0;
wire v$G2_12996_out0;
wire v$G2_12997_out0;
wire v$G2_12998_out0;
wire v$G2_12999_out0;
wire v$G2_13000_out0;
wire v$G2_13001_out0;
wire v$G2_13002_out0;
wire v$G2_13003_out0;
wire v$G2_13004_out0;
wire v$G2_13005_out0;
wire v$G2_13006_out0;
wire v$G2_13007_out0;
wire v$G2_13008_out0;
wire v$G2_13009_out0;
wire v$G2_13010_out0;
wire v$G2_13011_out0;
wire v$G2_13012_out0;
wire v$G2_13013_out0;
wire v$G2_13014_out0;
wire v$G2_13015_out0;
wire v$G2_13016_out0;
wire v$G2_13017_out0;
wire v$G2_13018_out0;
wire v$G2_13019_out0;
wire v$G2_13020_out0;
wire v$G2_13021_out0;
wire v$G2_13022_out0;
wire v$G2_13023_out0;
wire v$G2_13024_out0;
wire v$G2_13025_out0;
wire v$G2_13026_out0;
wire v$G2_13027_out0;
wire v$G2_13028_out0;
wire v$G2_13029_out0;
wire v$G2_13030_out0;
wire v$G2_13031_out0;
wire v$G2_13032_out0;
wire v$G2_13033_out0;
wire v$G2_13034_out0;
wire v$G2_13035_out0;
wire v$G2_13036_out0;
wire v$G2_13037_out0;
wire v$G2_13038_out0;
wire v$G2_13039_out0;
wire v$G2_13040_out0;
wire v$G2_13041_out0;
wire v$G2_13042_out0;
wire v$G2_13043_out0;
wire v$G2_13044_out0;
wire v$G2_13045_out0;
wire v$G2_13046_out0;
wire v$G2_13047_out0;
wire v$G2_13048_out0;
wire v$G2_13049_out0;
wire v$G2_13050_out0;
wire v$G2_13051_out0;
wire v$G2_13052_out0;
wire v$G2_13053_out0;
wire v$G2_13054_out0;
wire v$G2_13055_out0;
wire v$G2_13056_out0;
wire v$G2_13057_out0;
wire v$G2_13058_out0;
wire v$G2_13059_out0;
wire v$G2_13060_out0;
wire v$G2_13061_out0;
wire v$G2_13062_out0;
wire v$G2_13063_out0;
wire v$G2_13064_out0;
wire v$G2_13065_out0;
wire v$G2_13066_out0;
wire v$G2_13067_out0;
wire v$G2_13068_out0;
wire v$G2_13069_out0;
wire v$G2_13070_out0;
wire v$G2_13071_out0;
wire v$G2_13072_out0;
wire v$G2_13073_out0;
wire v$G2_13074_out0;
wire v$G2_13075_out0;
wire v$G2_13076_out0;
wire v$G2_13077_out0;
wire v$G2_13078_out0;
wire v$G2_13079_out0;
wire v$G2_13080_out0;
wire v$G2_13081_out0;
wire v$G2_13082_out0;
wire v$G2_13083_out0;
wire v$G2_13084_out0;
wire v$G2_13085_out0;
wire v$G2_13086_out0;
wire v$G2_13087_out0;
wire v$G2_13088_out0;
wire v$G2_13089_out0;
wire v$G2_13090_out0;
wire v$G2_13091_out0;
wire v$G2_13092_out0;
wire v$G2_13093_out0;
wire v$G2_13094_out0;
wire v$G2_13095_out0;
wire v$G2_13096_out0;
wire v$G2_13097_out0;
wire v$G2_13098_out0;
wire v$G2_13099_out0;
wire v$G2_13100_out0;
wire v$G2_13101_out0;
wire v$G2_13102_out0;
wire v$G2_13103_out0;
wire v$G2_13104_out0;
wire v$G2_13105_out0;
wire v$G2_13106_out0;
wire v$G2_13107_out0;
wire v$G2_13108_out0;
wire v$G2_13109_out0;
wire v$G2_13110_out0;
wire v$G2_13111_out0;
wire v$G2_13112_out0;
wire v$G2_13113_out0;
wire v$G2_13114_out0;
wire v$G2_13115_out0;
wire v$G2_13116_out0;
wire v$G2_13117_out0;
wire v$G2_13118_out0;
wire v$G2_13119_out0;
wire v$G2_13120_out0;
wire v$G2_13121_out0;
wire v$G2_13122_out0;
wire v$G2_13123_out0;
wire v$G2_13124_out0;
wire v$G2_13125_out0;
wire v$G2_13126_out0;
wire v$G2_13127_out0;
wire v$G2_13128_out0;
wire v$G2_13129_out0;
wire v$G2_13130_out0;
wire v$G2_13131_out0;
wire v$G2_13132_out0;
wire v$G2_13133_out0;
wire v$G2_13134_out0;
wire v$G2_13135_out0;
wire v$G2_13136_out0;
wire v$G2_13137_out0;
wire v$G2_13138_out0;
wire v$G2_13139_out0;
wire v$G2_13140_out0;
wire v$G2_13141_out0;
wire v$G2_13142_out0;
wire v$G2_13143_out0;
wire v$G2_13144_out0;
wire v$G2_13145_out0;
wire v$G2_13146_out0;
wire v$G2_13147_out0;
wire v$G2_13148_out0;
wire v$G2_13149_out0;
wire v$G2_13150_out0;
wire v$G2_13151_out0;
wire v$G2_13152_out0;
wire v$G2_13153_out0;
wire v$G2_13154_out0;
wire v$G2_13155_out0;
wire v$G2_13156_out0;
wire v$G2_13157_out0;
wire v$G2_13158_out0;
wire v$G2_13159_out0;
wire v$G2_13160_out0;
wire v$G2_13161_out0;
wire v$G2_13162_out0;
wire v$G2_13163_out0;
wire v$G2_13164_out0;
wire v$G2_13165_out0;
wire v$G2_13166_out0;
wire v$G2_13167_out0;
wire v$G2_13168_out0;
wire v$G2_13169_out0;
wire v$G2_13170_out0;
wire v$G2_13171_out0;
wire v$G2_13172_out0;
wire v$G2_13173_out0;
wire v$G2_13174_out0;
wire v$G2_13175_out0;
wire v$G2_13176_out0;
wire v$G2_13177_out0;
wire v$G2_13178_out0;
wire v$G2_13179_out0;
wire v$G2_13180_out0;
wire v$G2_13645_out0;
wire v$G2_13646_out0;
wire v$G2_1809_out0;
wire v$G2_1810_out0;
wire v$G2_1811_out0;
wire v$G2_1812_out0;
wire v$G2_1887_out0;
wire v$G2_1888_out0;
wire v$G2_2652_out0;
wire v$G2_2653_out0;
wire v$G2_2891_out0;
wire v$G2_2892_out0;
wire v$G2_2975_out0;
wire v$G2_2976_out0;
wire v$G2_2977_out0;
wire v$G2_2978_out0;
wire v$G2_3214_out0;
wire v$G2_3221_out0;
wire v$G2_3239_out0;
wire v$G2_3240_out0;
wire v$G2_3245_out0;
wire v$G2_3246_out0;
wire v$G2_4467_out0;
wire v$G2_4468_out0;
wire v$G2_4620_out0;
wire v$G2_4621_out0;
wire v$G2_4622_out0;
wire v$G2_4623_out0;
wire v$G2_4624_out0;
wire v$G2_4625_out0;
wire v$G2_4626_out0;
wire v$G2_4627_out0;
wire v$G2_4628_out0;
wire v$G2_4629_out0;
wire v$G2_4630_out0;
wire v$G2_4631_out0;
wire v$G2_4632_out0;
wire v$G2_4633_out0;
wire v$G2_4634_out0;
wire v$G2_4635_out0;
wire v$G2_4636_out0;
wire v$G2_4637_out0;
wire v$G2_4638_out0;
wire v$G2_4639_out0;
wire v$G2_4640_out0;
wire v$G2_4641_out0;
wire v$G2_4642_out0;
wire v$G2_4643_out0;
wire v$G2_4644_out0;
wire v$G2_4645_out0;
wire v$G2_4646_out0;
wire v$G2_4647_out0;
wire v$G2_4648_out0;
wire v$G2_4649_out0;
wire v$G2_5840_out0;
wire v$G2_5841_out0;
wire v$G2_6791_out0;
wire v$G2_6792_out0;
wire v$G2_6884_out0;
wire v$G2_6885_out0;
wire v$G2_7015_out0;
wire v$G2_7016_out0;
wire v$G2_7025_out0;
wire v$G2_7026_out0;
wire v$G2_7027_out0;
wire v$G2_7028_out0;
wire v$G30_183_out0;
wire v$G30_184_out0;
wire v$G35_10360_out0;
wire v$G35_10361_out0;
wire v$G35_10362_out0;
wire v$G35_10363_out0;
wire v$G36_3135_out0;
wire v$G36_3136_out0;
wire v$G36_3137_out0;
wire v$G36_3138_out0;
wire v$G37_6900_out0;
wire v$G37_6901_out0;
wire v$G37_6902_out0;
wire v$G37_6903_out0;
wire v$G38_3903_out0;
wire v$G38_3904_out0;
wire v$G38_3905_out0;
wire v$G38_3906_out0;
wire v$G3_10462_out0;
wire v$G3_13507_out0;
wire v$G3_13641_out0;
wire v$G3_13642_out0;
wire v$G3_1720_out0;
wire v$G3_1721_out0;
wire v$G3_17_out0;
wire v$G3_18_out0;
wire v$G3_1949_out0;
wire v$G3_1950_out0;
wire v$G3_206_out0;
wire v$G3_207_out0;
wire v$G3_208_out0;
wire v$G3_209_out0;
wire v$G3_241_out0;
wire v$G3_242_out0;
wire v$G3_243_out0;
wire v$G3_244_out0;
wire v$G3_245_out0;
wire v$G3_246_out0;
wire v$G3_247_out0;
wire v$G3_248_out0;
wire v$G3_249_out0;
wire v$G3_250_out0;
wire v$G3_251_out0;
wire v$G3_252_out0;
wire v$G3_253_out0;
wire v$G3_254_out0;
wire v$G3_255_out0;
wire v$G3_256_out0;
wire v$G3_257_out0;
wire v$G3_258_out0;
wire v$G3_259_out0;
wire v$G3_260_out0;
wire v$G3_261_out0;
wire v$G3_2621_out0;
wire v$G3_2622_out0;
wire v$G3_262_out0;
wire v$G3_263_out0;
wire v$G3_264_out0;
wire v$G3_265_out0;
wire v$G3_266_out0;
wire v$G3_267_out0;
wire v$G3_268_out0;
wire v$G3_2690_out0;
wire v$G3_2691_out0;
wire v$G3_269_out0;
wire v$G3_270_out0;
wire v$G3_2903_out0;
wire v$G3_2904_out0;
wire v$G3_2941_out0;
wire v$G3_2942_out0;
wire v$G3_3343_out0;
wire v$G3_3812_out0;
wire v$G3_3813_out0;
wire v$G3_3948_out0;
wire v$G3_3959_out0;
wire v$G3_3960_out0;
wire v$G3_6894_out0;
wire v$G3_6895_out0;
wire v$G3_6896_out0;
wire v$G3_6897_out0;
wire v$G3_7087_out0;
wire v$G3_7088_out0;
wire v$G3_7089_out0;
wire v$G3_7090_out0;
wire v$G3_8665_out0;
wire v$G3_8666_out0;
wire v$G4_10283_out0;
wire v$G4_10284_out0;
wire v$G4_10997_out0;
wire v$G4_10998_out0;
wire v$G4_10999_out0;
wire v$G4_11000_out0;
wire v$G4_12238_out0;
wire v$G4_12239_out0;
wire v$G4_12243_out0;
wire v$G4_12244_out0;
wire v$G4_13702_out0;
wire v$G4_13703_out0;
wire v$G4_1667_out0;
wire v$G4_1668_out0;
wire v$G4_1960_out0;
wire v$G4_1961_out0;
wire v$G4_1962_out0;
wire v$G4_1963_out0;
wire v$G4_219_out0;
wire v$G4_220_out0;
wire v$G4_2767_out0;
wire v$G4_2768_out0;
wire v$G4_2769_out0;
wire v$G4_2770_out0;
wire v$G4_3235_out0;
wire v$G4_3236_out0;
wire v$G4_341_out0;
wire v$G4_342_out0;
wire v$G4_343_out0;
wire v$G4_344_out0;
wire v$G4_345_out0;
wire v$G4_346_out0;
wire v$G4_347_out0;
wire v$G4_348_out0;
wire v$G4_349_out0;
wire v$G4_350_out0;
wire v$G4_351_out0;
wire v$G4_352_out0;
wire v$G4_353_out0;
wire v$G4_354_out0;
wire v$G4_355_out0;
wire v$G4_356_out0;
wire v$G4_357_out0;
wire v$G4_358_out0;
wire v$G4_359_out0;
wire v$G4_360_out0;
wire v$G4_361_out0;
wire v$G4_362_out0;
wire v$G4_363_out0;
wire v$G4_364_out0;
wire v$G4_365_out0;
wire v$G4_366_out0;
wire v$G4_367_out0;
wire v$G4_368_out0;
wire v$G4_369_out0;
wire v$G4_370_out0;
wire v$G4_381_out0;
wire v$G4_382_out0;
wire v$G4_4738_out0;
wire v$G4_4739_out0;
wire v$G4_4846_out0;
wire v$G4_4847_out0;
wire v$G4_6914_out0;
wire v$G4_6915_out0;
wire v$G5_10441_out0;
wire v$G5_10442_out0;
wire v$G5_10533_out0;
wire v$G5_10534_out0;
wire v$G5_10568_out0;
wire v$G5_10569_out0;
wire v$G5_10570_out0;
wire v$G5_10571_out0;
wire v$G5_10621_out0;
wire v$G5_10622_out0;
wire v$G5_10623_out0;
wire v$G5_10624_out0;
wire v$G5_10625_out0;
wire v$G5_10626_out0;
wire v$G5_10627_out0;
wire v$G5_10628_out0;
wire v$G5_10629_out0;
wire v$G5_10630_out0;
wire v$G5_10631_out0;
wire v$G5_10632_out0;
wire v$G5_10633_out0;
wire v$G5_10634_out0;
wire v$G5_10635_out0;
wire v$G5_10636_out0;
wire v$G5_10637_out0;
wire v$G5_10638_out0;
wire v$G5_10639_out0;
wire v$G5_10640_out0;
wire v$G5_10641_out0;
wire v$G5_10642_out0;
wire v$G5_10643_out0;
wire v$G5_10644_out0;
wire v$G5_10645_out0;
wire v$G5_10646_out0;
wire v$G5_10647_out0;
wire v$G5_10648_out0;
wire v$G5_10649_out0;
wire v$G5_10650_out0;
wire v$G5_10801_out0;
wire v$G5_10914_out0;
wire v$G5_10915_out0;
wire v$G5_10989_out0;
wire v$G5_1198_out0;
wire v$G5_229_out0;
wire v$G5_230_out0;
wire v$G5_2584_out0;
wire v$G5_2585_out0;
wire v$G5_2586_out0;
wire v$G5_2587_out0;
wire v$G5_2756_out0;
wire v$G5_2757_out0;
wire v$G5_2783_out0;
wire v$G5_2784_out0;
wire v$G5_2785_out0;
wire v$G5_2786_out0;
wire v$G5_4477_out0;
wire v$G5_4478_out0;
wire v$G5_454_out0;
wire v$G5_455_out0;
wire v$G5_638_out0;
wire v$G5_639_out0;
wire v$G5_7106_out0;
wire v$G5_7107_out0;
wire v$G6_11143_out0;
wire v$G6_11144_out0;
wire v$G6_1159_out0;
wire v$G6_1160_out0;
wire v$G6_1161_out0;
wire v$G6_1162_out0;
wire v$G6_13258_out0;
wire v$G6_13259_out0;
wire v$G6_13637_out0;
wire v$G6_13638_out0;
wire v$G6_13639_out0;
wire v$G6_13640_out0;
wire v$G6_2116_out0;
wire v$G6_2117_out0;
wire v$G6_2118_out0;
wire v$G6_2119_out0;
wire v$G6_2120_out0;
wire v$G6_2121_out0;
wire v$G6_2122_out0;
wire v$G6_2123_out0;
wire v$G6_2124_out0;
wire v$G6_2125_out0;
wire v$G6_2126_out0;
wire v$G6_2127_out0;
wire v$G6_2128_out0;
wire v$G6_2129_out0;
wire v$G6_2130_out0;
wire v$G6_2131_out0;
wire v$G6_2132_out0;
wire v$G6_2133_out0;
wire v$G6_2134_out0;
wire v$G6_2135_out0;
wire v$G6_2136_out0;
wire v$G6_2137_out0;
wire v$G6_2138_out0;
wire v$G6_2139_out0;
wire v$G6_2140_out0;
wire v$G6_2141_out0;
wire v$G6_2142_out0;
wire v$G6_2143_out0;
wire v$G6_2144_out0;
wire v$G6_2145_out0;
wire v$G6_2416_out0;
wire v$G6_2417_out0;
wire v$G6_2905_out0;
wire v$G6_2906_out0;
wire v$G6_327_out0;
wire v$G6_328_out0;
wire v$G6_4531_out0;
wire v$G6_4818_out0;
wire v$G6_8834_out0;
wire v$G6_8835_out0;
wire v$G6_8836_out0;
wire v$G6_8837_out0;
wire v$G7_10332_out0;
wire v$G7_11095_out0;
wire v$G7_11262_out0;
wire v$G7_11263_out0;
wire v$G7_11264_out0;
wire v$G7_11265_out0;
wire v$G7_11266_out0;
wire v$G7_11267_out0;
wire v$G7_11268_out0;
wire v$G7_11269_out0;
wire v$G7_11270_out0;
wire v$G7_11271_out0;
wire v$G7_11272_out0;
wire v$G7_11273_out0;
wire v$G7_11274_out0;
wire v$G7_11275_out0;
wire v$G7_11276_out0;
wire v$G7_11277_out0;
wire v$G7_11278_out0;
wire v$G7_11279_out0;
wire v$G7_11280_out0;
wire v$G7_11281_out0;
wire v$G7_11282_out0;
wire v$G7_11283_out0;
wire v$G7_11284_out0;
wire v$G7_11285_out0;
wire v$G7_11286_out0;
wire v$G7_11287_out0;
wire v$G7_11288_out0;
wire v$G7_11289_out0;
wire v$G7_11290_out0;
wire v$G7_11291_out0;
wire v$G7_1197_out0;
wire v$G7_1684_out0;
wire v$G7_1685_out0;
wire v$G7_169_out0;
wire v$G7_170_out0;
wire v$G7_2455_out0;
wire v$G7_2779_out0;
wire v$G7_2780_out0;
wire v$G7_2781_out0;
wire v$G7_2782_out0;
wire v$G7_4474_out0;
wire v$G7_4475_out0;
wire v$G7_4821_out0;
wire v$G7_4822_out0;
wire v$G7_6862_out0;
wire v$G7_6863_out0;
wire v$G7_8655_out0;
wire v$G7_8656_out0;
wire v$G7_8657_out0;
wire v$G7_8658_out0;
wire v$G8_10609_out0;
wire v$G8_10610_out0;
wire v$G8_10611_out0;
wire v$G8_10612_out0;
wire v$G8_10769_out0;
wire v$G8_10770_out0;
wire v$G8_1215_out0;
wire v$G8_1216_out0;
wire v$G8_1217_out0;
wire v$G8_1218_out0;
wire v$G8_16_out0;
wire v$G8_1765_out0;
wire v$G8_1766_out0;
wire v$G8_2024_out0;
wire v$G8_2025_out0;
wire v$G8_2472_out0;
wire v$G8_2473_out0;
wire v$G8_2474_out0;
wire v$G8_2475_out0;
wire v$G8_2476_out0;
wire v$G8_2477_out0;
wire v$G8_2478_out0;
wire v$G8_2479_out0;
wire v$G8_2480_out0;
wire v$G8_2481_out0;
wire v$G8_2482_out0;
wire v$G8_2483_out0;
wire v$G8_2484_out0;
wire v$G8_2485_out0;
wire v$G8_2486_out0;
wire v$G8_2487_out0;
wire v$G8_2488_out0;
wire v$G8_2489_out0;
wire v$G8_2490_out0;
wire v$G8_2491_out0;
wire v$G8_2492_out0;
wire v$G8_2493_out0;
wire v$G8_2494_out0;
wire v$G8_2495_out0;
wire v$G8_2496_out0;
wire v$G8_2497_out0;
wire v$G8_2498_out0;
wire v$G8_2499_out0;
wire v$G8_2500_out0;
wire v$G8_2501_out0;
wire v$G8_2623_out0;
wire v$G8_2624_out0;
wire v$G8_2644_out0;
wire v$G8_4453_out0;
wire v$G8_4454_out0;
wire v$G8_548_out0;
wire v$G8_549_out0;
wire v$G8_550_out0;
wire v$G8_551_out0;
wire v$G8_7103_out0;
wire v$G9_10291_out0;
wire v$G9_10292_out0;
wire v$G9_10293_out0;
wire v$G9_10294_out0;
wire v$G9_10572_out0;
wire v$G9_10573_out0;
wire v$G9_10574_out0;
wire v$G9_10575_out0;
wire v$G9_10576_out0;
wire v$G9_10577_out0;
wire v$G9_10578_out0;
wire v$G9_10579_out0;
wire v$G9_10580_out0;
wire v$G9_10581_out0;
wire v$G9_10582_out0;
wire v$G9_10583_out0;
wire v$G9_10584_out0;
wire v$G9_10585_out0;
wire v$G9_10586_out0;
wire v$G9_10587_out0;
wire v$G9_10588_out0;
wire v$G9_10589_out0;
wire v$G9_10590_out0;
wire v$G9_10591_out0;
wire v$G9_10592_out0;
wire v$G9_10593_out0;
wire v$G9_10594_out0;
wire v$G9_10595_out0;
wire v$G9_10596_out0;
wire v$G9_10597_out0;
wire v$G9_10598_out0;
wire v$G9_10599_out0;
wire v$G9_10600_out0;
wire v$G9_10601_out0;
wire v$G9_13285_out0;
wire v$G9_13286_out0;
wire v$G9_13287_out0;
wire v$G9_13288_out0;
wire v$G9_13340_out0;
wire v$G9_13341_out0;
wire v$G9_13564_out0;
wire v$G9_13655_out0;
wire v$G9_1671_out0;
wire v$G9_1672_out0;
wire v$G9_223_out0;
wire v$G9_2332_out0;
wire v$G9_2333_out0;
wire v$G9_2895_out0;
wire v$G9_2896_out0;
wire v$G9_2897_out0;
wire v$G9_2898_out0;
wire v$G9_407_out0;
wire v$G9_408_out0;
wire v$G9_411_out0;
wire v$G9_412_out0;
wire v$IN_2466_out0;
wire v$IR15_2464_out0;
wire v$IR15_2465_out0;
wire v$JEQZ_10514_out0;
wire v$JEQZ_10515_out0;
wire v$JEQZ_2981_out0;
wire v$JEQZ_2982_out0;
wire v$JEQ_10496_out0;
wire v$JEQ_10497_out0;
wire v$JEQ_13560_out0;
wire v$JEQ_13561_out0;
wire v$JEQ_2234_out0;
wire v$JEQ_2235_out0;
wire v$JEQ_4445_out0;
wire v$JEQ_4446_out0;
wire v$JEQ_8806_out0;
wire v$JEQ_8807_out0;
wire v$JMIN_1205_out0;
wire v$JMIN_1206_out0;
wire v$JMIN_2662_out0;
wire v$JMIN_2663_out0;
wire v$JMI_13349_out0;
wire v$JMI_13350_out0;
wire v$JMI_1939_out0;
wire v$JMI_1940_out0;
wire v$JMI_3212_out0;
wire v$JMI_3213_out0;
wire v$JMI_8679_out0;
wire v$JMI_8680_out0;
wire v$JMI_88_out0;
wire v$JMI_89_out0;
wire v$JMP_2668_out0;
wire v$JMP_2669_out0;
wire v$JMP_3233_out0;
wire v$JMP_3234_out0;
wire v$JMP_546_out0;
wire v$JMP_547_out0;
wire v$JMP_7077_out0;
wire v$JMP_7078_out0;
wire v$JMP_8825_out0;
wire v$JMP_8826_out0;
wire v$JUMP_2187_out0;
wire v$JUMP_2188_out0;
wire v$LDR$STR0_10349_out0;
wire v$LDR$STR1_13616_out0;
wire v$LOAD_231_out0;
wire v$LOAD_232_out0;
wire v$LOAD_2899_out0;
wire v$LOAD_2900_out0;
wire v$LOAD_3115_out0;
wire v$LOAD_3116_out0;
wire v$LOAD_3949_out0;
wire v$LOAD_3950_out0;
wire v$LOAD_7110_out0;
wire v$LOAD_7111_out0;
wire v$LOAD_8765_out0;
wire v$LOAD_8766_out0;
wire v$LS0_4548_out0;
wire v$LS1_3169_out0;
wire v$LSL_1861_out0;
wire v$LSL_1862_out0;
wire v$LSL_2842_out0;
wire v$LSL_2843_out0;
wire v$LSL_3047_out0;
wire v$LSL_3048_out0;
wire v$LSL_3182_out0;
wire v$LSL_3183_out0;
wire v$LSR_1174_out0;
wire v$LSR_1175_out0;
wire v$LSR_13331_out0;
wire v$LSR_13332_out0;
wire v$LSR_418_out0;
wire v$LSR_419_out0;
wire v$LSR_6912_out0;
wire v$LSR_6913_out0;
wire v$LS_1202_out0;
wire v$LS_1203_out0;
wire v$LS_202_out0;
wire v$LS_203_out0;
wire v$LS_204_out0;
wire v$LS_205_out0;
wire v$LS_2864_out0;
wire v$LS_2865_out0;
wire v$MI_10833_out0;
wire v$MI_10834_out0;
wire v$MI_2612_out0;
wire v$MI_2613_out0;
wire v$MI_560_out0;
wire v$MI_561_out0;
wire v$MOV_10389_out0;
wire v$MOV_10390_out0;
wire v$MOV_196_out0;
wire v$MOV_197_out0;
wire v$MULTI$INSTRUCTION_13308_out0;
wire v$MULTI$INSTRUCTION_13309_out0;
wire v$MULTI$INSTRUCTION_13323_out0;
wire v$MULTI$INSTRUCTION_13324_out0;
wire v$MULTI$INSTRUCTION_2451_out0;
wire v$MULTI$INSTRUCTION_2452_out0;
wire v$MULTI$INSTRUCTION_3953_out0;
wire v$MULTI$INSTRUCTION_3954_out0;
wire v$MULTI$INSTRUCTION_619_out0;
wire v$MULTI$INSTRUCTION_620_out0;
wire v$MULTI$OPCODE_10797_out0;
wire v$MULTI$OPCODE_10798_out0;
wire v$MULTI$OPCODE_11096_out0;
wire v$MULTI$OPCODE_11097_out0;
wire v$MULTI$OPCODE_3020_out0;
wire v$MULTI$OPCODE_3021_out0;
wire v$MUX$ENABLE_2349_out0;
wire v$MUX1_2625_out0;
wire v$MUX1_650_out0;
wire v$MUX2_1180_out0;
wire v$MUX2_4448_out0;
wire v$MUX3_10994_out0;
wire v$MUX3_7140_out0;
wire v$MUX3_8817_out0;
wire v$MUX3_8818_out0;
wire v$MUX4_3219_out0;
wire v$MUX5_10260_out0;
wire v$MUX5_10261_out0;
wire v$MUX5_13348_out0;
wire v$MUX5_7678_out0;
wire v$MUX6_10976_out0;
wire v$MUX6_8757_out0;
wire v$MUX6_8758_out0;
wire v$MUX7_10448_out0;
wire v$MUX8_2697_out0;
wire v$MUX9_166_out0;
wire v$NEGATIVE_11256_out0;
wire v$NEGATIVE_11257_out0;
wire v$NORMAL0_2307_out0;
wire v$NORMAL1_6790_out0;
wire v$NORMAL_10256_out0;
wire v$NORMAL_10257_out0;
wire v$NORMAL_13429_out0;
wire v$NORMAL_13430_out0;
wire v$NORMAL_181_out0;
wire v$NORMAL_182_out0;
wire v$NORMAL_3353_out0;
wire v$NORMAL_3354_out0;
wire v$NORMAL_7114_out0;
wire v$NORMAL_7115_out0;
wire v$NOTUSED1_10684_out0;
wire v$NOTUSED1_10685_out0;
wire v$NOTUSED2_5794_out0;
wire v$NOTUSED2_5795_out0;
wire v$NOTUSED3_10550_out0;
wire v$NOTUSED3_10551_out0;
wire v$NOTUSED4_10530_out0;
wire v$NOTUSED4_10531_out0;
wire v$NOTUSED_10835_out0;
wire v$NOTUSED_10836_out0;
wire v$NOTUSED_1968_out0;
wire v$NOTUSED_1969_out0;
wire v$NOTUSED_325_out0;
wire v$NOTUSED_326_out0;
wire v$NOTUSED_4463_out0;
wire v$NOTUSED_4464_out0;
wire v$NOTUSED_4609_out0;
wire v$OP2$SIGN_10839_out0;
wire v$OP2$SIGN_10840_out0;
wire v$OP2$SIGN_11208_out0;
wire v$OP2$SIGN_11209_out0;
wire v$OUTSTREAM_2097_out0;
wire v$OUT_22_out0;
wire v$OVERFLOW_10492_out0;
wire v$OVERFLOW_10493_out0;
wire v$P_10682_out0;
wire v$P_10683_out0;
wire v$Q0_11198_out0;
wire v$Q0_11199_out0;
wire v$Q0_11200_out0;
wire v$Q0_11201_out0;
wire v$Q0_13351_out0;
wire v$Q0_4470_out0;
wire v$Q0_4471_out0;
wire v$Q0_4472_out0;
wire v$Q0_4473_out0;
wire v$Q0_625_out0;
wire v$Q0_626_out0;
wire v$Q1_2112_out0;
wire v$Q1_307_out0;
wire v$Q1_308_out0;
wire v$Q1_3993_out0;
wire v$Q1_6906_out0;
wire v$Q1_6907_out0;
wire v$Q1_6908_out0;
wire v$Q1_6909_out0;
wire v$Q1_8859_out0;
wire v$Q1_8860_out0;
wire v$Q1_8861_out0;
wire v$Q1_8862_out0;
wire v$Q2_1676_out0;
wire v$Q2_1677_out0;
wire v$Q2_1678_out0;
wire v$Q2_1679_out0;
wire v$Q2_6880_out0;
wire v$Q2_6881_out0;
wire v$Q2_6882_out0;
wire v$Q2_6883_out0;
wire v$Q3_10518_out0;
wire v$Q3_10519_out0;
wire v$Q3_10520_out0;
wire v$Q3_10521_out0;
wire v$Q3_8737_out0;
wire v$Q3_8738_out0;
wire v$Q3_8739_out0;
wire v$Q3_8740_out0;
wire v$Q6_1889_out0;
wire v$Q6_1890_out0;
wire v$Q6_1891_out0;
wire v$Q6_1892_out0;
wire v$Q7_6888_out0;
wire v$Q7_6889_out0;
wire v$Q7_6890_out0;
wire v$Q7_6891_out0;
wire v$Q_291_out0;
wire v$Q_292_out0;
wire v$Q_293_out0;
wire v$Q_294_out0;
wire v$Q_295_out0;
wire v$Q_296_out0;
wire v$Q_297_out0;
wire v$Q_298_out0;
wire v$Q_299_out0;
wire v$Q_300_out0;
wire v$Q_301_out0;
wire v$Q_302_out0;
wire v$Q_303_out0;
wire v$Q_304_out0;
wire v$Q_305_out0;
wire v$Q_306_out0;
wire v$RAMWEN_10701_out0;
wire v$RAMWEN_10702_out0;
wire v$RD$SIGN_2405_out0;
wire v$RD$SIGN_2406_out0;
wire v$RD$SIGN_285_out0;
wire v$RD$SIGN_286_out0;
wire v$RDN_3349_out0;
wire v$RDN_3351_out0;
wire v$RDN_4496_out0;
wire v$RDN_4497_out0;
wire v$RDN_4498_out0;
wire v$RDN_4499_out0;
wire v$RDN_4500_out0;
wire v$RDN_4501_out0;
wire v$RDN_4502_out0;
wire v$RDN_4503_out0;
wire v$RDN_4504_out0;
wire v$RDN_4505_out0;
wire v$RDN_4506_out0;
wire v$RDN_4507_out0;
wire v$RDN_4508_out0;
wire v$RDN_4509_out0;
wire v$RDN_4510_out0;
wire v$RDN_4511_out0;
wire v$RDN_4512_out0;
wire v$RDN_4513_out0;
wire v$RDN_4514_out0;
wire v$RDN_4515_out0;
wire v$RDN_4516_out0;
wire v$RDN_4517_out0;
wire v$RDN_4518_out0;
wire v$RDN_4519_out0;
wire v$RDN_4520_out0;
wire v$RDN_4521_out0;
wire v$RDN_4522_out0;
wire v$RDN_4523_out0;
wire v$RDN_4524_out0;
wire v$RDN_4525_out0;
wire v$RD_13567_out0;
wire v$RD_13568_out0;
wire v$RD_13569_out0;
wire v$RD_13570_out0;
wire v$RD_13571_out0;
wire v$RD_13572_out0;
wire v$RD_13573_out0;
wire v$RD_13574_out0;
wire v$RD_13575_out0;
wire v$RD_13576_out0;
wire v$RD_13577_out0;
wire v$RD_13578_out0;
wire v$RD_13579_out0;
wire v$RD_13580_out0;
wire v$RD_13581_out0;
wire v$RD_13582_out0;
wire v$RD_13583_out0;
wire v$RD_13584_out0;
wire v$RD_13585_out0;
wire v$RD_13586_out0;
wire v$RD_13587_out0;
wire v$RD_13588_out0;
wire v$RD_13589_out0;
wire v$RD_13590_out0;
wire v$RD_13591_out0;
wire v$RD_13592_out0;
wire v$RD_13593_out0;
wire v$RD_13594_out0;
wire v$RD_13595_out0;
wire v$RD_13596_out0;
wire v$RD_5862_out0;
wire v$RD_5863_out0;
wire v$RD_5864_out0;
wire v$RD_5865_out0;
wire v$RD_5866_out0;
wire v$RD_5867_out0;
wire v$RD_5868_out0;
wire v$RD_5869_out0;
wire v$RD_5870_out0;
wire v$RD_5871_out0;
wire v$RD_5872_out0;
wire v$RD_5873_out0;
wire v$RD_5874_out0;
wire v$RD_5875_out0;
wire v$RD_5876_out0;
wire v$RD_5877_out0;
wire v$RD_5878_out0;
wire v$RD_5879_out0;
wire v$RD_5880_out0;
wire v$RD_5881_out0;
wire v$RD_5882_out0;
wire v$RD_5883_out0;
wire v$RD_5884_out0;
wire v$RD_5885_out0;
wire v$RD_5886_out0;
wire v$RD_5887_out0;
wire v$RD_5888_out0;
wire v$RD_5889_out0;
wire v$RD_5890_out0;
wire v$RD_5891_out0;
wire v$RD_5892_out0;
wire v$RD_5893_out0;
wire v$RD_5894_out0;
wire v$RD_5895_out0;
wire v$RD_5896_out0;
wire v$RD_5897_out0;
wire v$RD_5898_out0;
wire v$RD_5899_out0;
wire v$RD_5900_out0;
wire v$RD_5901_out0;
wire v$RD_5902_out0;
wire v$RD_5903_out0;
wire v$RD_5904_out0;
wire v$RD_5905_out0;
wire v$RD_5906_out0;
wire v$RD_5907_out0;
wire v$RD_5908_out0;
wire v$RD_5909_out0;
wire v$RD_5910_out0;
wire v$RD_5911_out0;
wire v$RD_5912_out0;
wire v$RD_5913_out0;
wire v$RD_5914_out0;
wire v$RD_5915_out0;
wire v$RD_5916_out0;
wire v$RD_5917_out0;
wire v$RD_5918_out0;
wire v$RD_5919_out0;
wire v$RD_5920_out0;
wire v$RD_5921_out0;
wire v$RD_5922_out0;
wire v$RD_5923_out0;
wire v$RD_5924_out0;
wire v$RD_5925_out0;
wire v$RD_5926_out0;
wire v$RD_5927_out0;
wire v$RD_5928_out0;
wire v$RD_5929_out0;
wire v$RD_5930_out0;
wire v$RD_5931_out0;
wire v$RD_5932_out0;
wire v$RD_5933_out0;
wire v$RD_5934_out0;
wire v$RD_5935_out0;
wire v$RD_5936_out0;
wire v$RD_5937_out0;
wire v$RD_5938_out0;
wire v$RD_5939_out0;
wire v$RD_5940_out0;
wire v$RD_5941_out0;
wire v$RD_5942_out0;
wire v$RD_5943_out0;
wire v$RD_5944_out0;
wire v$RD_5945_out0;
wire v$RD_5946_out0;
wire v$RD_5947_out0;
wire v$RD_5948_out0;
wire v$RD_5949_out0;
wire v$RD_5950_out0;
wire v$RD_5951_out0;
wire v$RD_5952_out0;
wire v$RD_5953_out0;
wire v$RD_5954_out0;
wire v$RD_5955_out0;
wire v$RD_5956_out0;
wire v$RD_5957_out0;
wire v$RD_5958_out0;
wire v$RD_5959_out0;
wire v$RD_5960_out0;
wire v$RD_5961_out0;
wire v$RD_5962_out0;
wire v$RD_5963_out0;
wire v$RD_5964_out0;
wire v$RD_5965_out0;
wire v$RD_5966_out0;
wire v$RD_5967_out0;
wire v$RD_5968_out0;
wire v$RD_5969_out0;
wire v$RD_5970_out0;
wire v$RD_5971_out0;
wire v$RD_5972_out0;
wire v$RD_5973_out0;
wire v$RD_5974_out0;
wire v$RD_5975_out0;
wire v$RD_5976_out0;
wire v$RD_5977_out0;
wire v$RD_5978_out0;
wire v$RD_5979_out0;
wire v$RD_5980_out0;
wire v$RD_5981_out0;
wire v$RD_5982_out0;
wire v$RD_5983_out0;
wire v$RD_5984_out0;
wire v$RD_5985_out0;
wire v$RD_5986_out0;
wire v$RD_5987_out0;
wire v$RD_5988_out0;
wire v$RD_5989_out0;
wire v$RD_5990_out0;
wire v$RD_5991_out0;
wire v$RD_5992_out0;
wire v$RD_5993_out0;
wire v$RD_5994_out0;
wire v$RD_5995_out0;
wire v$RD_5996_out0;
wire v$RD_5997_out0;
wire v$RD_5998_out0;
wire v$RD_5999_out0;
wire v$RD_6000_out0;
wire v$RD_6001_out0;
wire v$RD_6002_out0;
wire v$RD_6003_out0;
wire v$RD_6004_out0;
wire v$RD_6005_out0;
wire v$RD_6006_out0;
wire v$RD_6007_out0;
wire v$RD_6008_out0;
wire v$RD_6009_out0;
wire v$RD_6010_out0;
wire v$RD_6011_out0;
wire v$RD_6012_out0;
wire v$RD_6013_out0;
wire v$RD_6014_out0;
wire v$RD_6015_out0;
wire v$RD_6016_out0;
wire v$RD_6017_out0;
wire v$RD_6018_out0;
wire v$RD_6019_out0;
wire v$RD_6020_out0;
wire v$RD_6021_out0;
wire v$RD_6022_out0;
wire v$RD_6023_out0;
wire v$RD_6024_out0;
wire v$RD_6025_out0;
wire v$RD_6026_out0;
wire v$RD_6027_out0;
wire v$RD_6028_out0;
wire v$RD_6029_out0;
wire v$RD_6030_out0;
wire v$RD_6031_out0;
wire v$RD_6032_out0;
wire v$RD_6033_out0;
wire v$RD_6034_out0;
wire v$RD_6035_out0;
wire v$RD_6036_out0;
wire v$RD_6037_out0;
wire v$RD_6038_out0;
wire v$RD_6039_out0;
wire v$RD_6040_out0;
wire v$RD_6041_out0;
wire v$RD_6042_out0;
wire v$RD_6043_out0;
wire v$RD_6044_out0;
wire v$RD_6045_out0;
wire v$RD_6046_out0;
wire v$RD_6047_out0;
wire v$RD_6048_out0;
wire v$RD_6049_out0;
wire v$RD_6050_out0;
wire v$RD_6051_out0;
wire v$RD_6052_out0;
wire v$RD_6053_out0;
wire v$RD_6054_out0;
wire v$RD_6055_out0;
wire v$RD_6056_out0;
wire v$RD_6057_out0;
wire v$RD_6058_out0;
wire v$RD_6059_out0;
wire v$RD_6060_out0;
wire v$RD_6061_out0;
wire v$RD_6062_out0;
wire v$RD_6063_out0;
wire v$RD_6064_out0;
wire v$RD_6065_out0;
wire v$RD_6066_out0;
wire v$RD_6067_out0;
wire v$RD_6068_out0;
wire v$RD_6069_out0;
wire v$RD_6070_out0;
wire v$RD_6071_out0;
wire v$RD_6072_out0;
wire v$RD_6073_out0;
wire v$RD_6074_out0;
wire v$RD_6075_out0;
wire v$RD_6076_out0;
wire v$RD_6077_out0;
wire v$RD_6078_out0;
wire v$RD_6079_out0;
wire v$RD_6080_out0;
wire v$RD_6081_out0;
wire v$RD_6082_out0;
wire v$RD_6083_out0;
wire v$RD_6084_out0;
wire v$RD_6085_out0;
wire v$RD_6086_out0;
wire v$RD_6087_out0;
wire v$RD_6088_out0;
wire v$RD_6089_out0;
wire v$RD_6090_out0;
wire v$RD_6091_out0;
wire v$RD_6092_out0;
wire v$RD_6093_out0;
wire v$RD_6094_out0;
wire v$RD_6095_out0;
wire v$RD_6096_out0;
wire v$RD_6097_out0;
wire v$RD_6098_out0;
wire v$RD_6099_out0;
wire v$RD_6100_out0;
wire v$RD_6101_out0;
wire v$RD_6102_out0;
wire v$RD_6103_out0;
wire v$RD_6104_out0;
wire v$RD_6105_out0;
wire v$RD_6106_out0;
wire v$RD_6107_out0;
wire v$RD_6108_out0;
wire v$RD_6109_out0;
wire v$RD_6110_out0;
wire v$RD_6111_out0;
wire v$RD_6112_out0;
wire v$RD_6113_out0;
wire v$RD_6114_out0;
wire v$RD_6115_out0;
wire v$RD_6116_out0;
wire v$RD_6117_out0;
wire v$RD_6118_out0;
wire v$RD_6119_out0;
wire v$RD_6120_out0;
wire v$RD_6121_out0;
wire v$RD_6122_out0;
wire v$RD_6123_out0;
wire v$RD_6124_out0;
wire v$RD_6125_out0;
wire v$RD_6126_out0;
wire v$RD_6127_out0;
wire v$RD_6128_out0;
wire v$RD_6129_out0;
wire v$RD_6130_out0;
wire v$RD_6131_out0;
wire v$RD_6132_out0;
wire v$RD_6133_out0;
wire v$RD_6134_out0;
wire v$RD_6135_out0;
wire v$RD_6136_out0;
wire v$RD_6137_out0;
wire v$RD_6138_out0;
wire v$RD_6139_out0;
wire v$RD_6140_out0;
wire v$RD_6141_out0;
wire v$RD_6142_out0;
wire v$RD_6143_out0;
wire v$RD_6144_out0;
wire v$RD_6145_out0;
wire v$RD_6146_out0;
wire v$RD_6147_out0;
wire v$RD_6148_out0;
wire v$RD_6149_out0;
wire v$RD_6150_out0;
wire v$RD_6151_out0;
wire v$RD_6152_out0;
wire v$RD_6153_out0;
wire v$RD_6154_out0;
wire v$RD_6155_out0;
wire v$RD_6156_out0;
wire v$RD_6157_out0;
wire v$RD_6158_out0;
wire v$RD_6159_out0;
wire v$RD_6160_out0;
wire v$RD_6161_out0;
wire v$RD_6162_out0;
wire v$RD_6163_out0;
wire v$RD_6164_out0;
wire v$RD_6165_out0;
wire v$RD_6166_out0;
wire v$RD_6167_out0;
wire v$RD_6168_out0;
wire v$RD_6169_out0;
wire v$RD_6170_out0;
wire v$RD_6171_out0;
wire v$RD_6172_out0;
wire v$RD_6173_out0;
wire v$RD_6174_out0;
wire v$RD_6175_out0;
wire v$RD_6176_out0;
wire v$RD_6177_out0;
wire v$RD_6178_out0;
wire v$RD_6179_out0;
wire v$RD_6180_out0;
wire v$RD_6181_out0;
wire v$RD_6182_out0;
wire v$RD_6183_out0;
wire v$RD_6184_out0;
wire v$RD_6185_out0;
wire v$RD_6186_out0;
wire v$RD_6187_out0;
wire v$RD_6188_out0;
wire v$RD_6189_out0;
wire v$RD_6190_out0;
wire v$RD_6191_out0;
wire v$RD_6192_out0;
wire v$RD_6193_out0;
wire v$RD_6194_out0;
wire v$RD_6195_out0;
wire v$RD_6196_out0;
wire v$RD_6197_out0;
wire v$RD_6198_out0;
wire v$RD_6199_out0;
wire v$RD_6200_out0;
wire v$RD_6201_out0;
wire v$RD_6202_out0;
wire v$RD_6203_out0;
wire v$RD_6204_out0;
wire v$RD_6205_out0;
wire v$RD_6206_out0;
wire v$RD_6207_out0;
wire v$RD_6208_out0;
wire v$RD_6209_out0;
wire v$RD_6210_out0;
wire v$RD_6211_out0;
wire v$RD_6212_out0;
wire v$RD_6213_out0;
wire v$RD_6214_out0;
wire v$RD_6215_out0;
wire v$RD_6216_out0;
wire v$RD_6217_out0;
wire v$RD_6218_out0;
wire v$RD_6219_out0;
wire v$RD_6220_out0;
wire v$RD_6221_out0;
wire v$RD_6222_out0;
wire v$RD_6223_out0;
wire v$RD_6224_out0;
wire v$RD_6225_out0;
wire v$RD_6226_out0;
wire v$RD_6227_out0;
wire v$RD_6228_out0;
wire v$RD_6229_out0;
wire v$RD_6230_out0;
wire v$RD_6231_out0;
wire v$RD_6232_out0;
wire v$RD_6233_out0;
wire v$RD_6234_out0;
wire v$RD_6235_out0;
wire v$RD_6236_out0;
wire v$RD_6237_out0;
wire v$RD_6238_out0;
wire v$RD_6239_out0;
wire v$RD_6240_out0;
wire v$RD_6241_out0;
wire v$RD_6242_out0;
wire v$RD_6243_out0;
wire v$RD_6244_out0;
wire v$RD_6245_out0;
wire v$RD_6246_out0;
wire v$RD_6247_out0;
wire v$RD_6248_out0;
wire v$RD_6249_out0;
wire v$RD_6250_out0;
wire v$RD_6251_out0;
wire v$RD_6252_out0;
wire v$RD_6253_out0;
wire v$RD_6254_out0;
wire v$RD_6255_out0;
wire v$RD_6256_out0;
wire v$RD_6257_out0;
wire v$RD_6258_out0;
wire v$RD_6259_out0;
wire v$RD_6260_out0;
wire v$RD_6261_out0;
wire v$RD_6262_out0;
wire v$RD_6263_out0;
wire v$RD_6264_out0;
wire v$RD_6265_out0;
wire v$RD_6266_out0;
wire v$RD_6267_out0;
wire v$RD_6268_out0;
wire v$RD_6269_out0;
wire v$RD_6270_out0;
wire v$RD_6271_out0;
wire v$RD_6272_out0;
wire v$RD_6273_out0;
wire v$RD_6274_out0;
wire v$RD_6275_out0;
wire v$RD_6276_out0;
wire v$RD_6277_out0;
wire v$RD_6278_out0;
wire v$RD_6279_out0;
wire v$RD_6280_out0;
wire v$RD_6281_out0;
wire v$RD_6282_out0;
wire v$RD_6283_out0;
wire v$RD_6284_out0;
wire v$RD_6285_out0;
wire v$RD_6286_out0;
wire v$RD_6287_out0;
wire v$RD_6288_out0;
wire v$RD_6289_out0;
wire v$RD_6290_out0;
wire v$RD_6291_out0;
wire v$RD_6292_out0;
wire v$RD_6293_out0;
wire v$RD_6294_out0;
wire v$RD_6295_out0;
wire v$RD_6296_out0;
wire v$RD_6297_out0;
wire v$RD_6298_out0;
wire v$RD_6299_out0;
wire v$RD_6300_out0;
wire v$RD_6301_out0;
wire v$RD_6302_out0;
wire v$RD_6303_out0;
wire v$RD_6304_out0;
wire v$RD_6305_out0;
wire v$RD_6306_out0;
wire v$RD_6307_out0;
wire v$RD_6308_out0;
wire v$RD_6309_out0;
wire v$RD_6310_out0;
wire v$RD_6311_out0;
wire v$RD_6312_out0;
wire v$RD_6313_out0;
wire v$RD_6314_out0;
wire v$RD_6315_out0;
wire v$RD_6316_out0;
wire v$RD_6317_out0;
wire v$RD_6318_out0;
wire v$RD_6319_out0;
wire v$RD_6320_out0;
wire v$RD_6321_out0;
wire v$RD_6322_out0;
wire v$RD_6323_out0;
wire v$RD_6324_out0;
wire v$RD_6325_out0;
wire v$RD_6326_out0;
wire v$RD_6327_out0;
wire v$RD_6328_out0;
wire v$RD_6329_out0;
wire v$RD_6330_out0;
wire v$RD_6331_out0;
wire v$RD_6332_out0;
wire v$RD_6333_out0;
wire v$RD_6334_out0;
wire v$RD_6335_out0;
wire v$RD_6336_out0;
wire v$RD_6337_out0;
wire v$RD_6338_out0;
wire v$RD_6339_out0;
wire v$RD_6340_out0;
wire v$RD_6341_out0;
wire v$RD_6342_out0;
wire v$RD_6343_out0;
wire v$RD_6344_out0;
wire v$RD_6345_out0;
wire v$RD_6346_out0;
wire v$RD_6347_out0;
wire v$RD_6348_out0;
wire v$RD_6349_out0;
wire v$RD_6350_out0;
wire v$RD_6351_out0;
wire v$RD_6352_out0;
wire v$RD_6353_out0;
wire v$RD_6354_out0;
wire v$RD_6355_out0;
wire v$RD_6356_out0;
wire v$RD_6357_out0;
wire v$RD_6358_out0;
wire v$RD_6359_out0;
wire v$RD_6360_out0;
wire v$RD_6361_out0;
wire v$RD_6362_out0;
wire v$RD_6363_out0;
wire v$RD_6364_out0;
wire v$RD_6365_out0;
wire v$RD_6366_out0;
wire v$RD_6367_out0;
wire v$RD_6368_out0;
wire v$RD_6369_out0;
wire v$RD_6370_out0;
wire v$RD_6371_out0;
wire v$RD_6372_out0;
wire v$RD_6373_out0;
wire v$RD_6374_out0;
wire v$RD_6375_out0;
wire v$RD_6376_out0;
wire v$RD_6377_out0;
wire v$RD_6378_out0;
wire v$RD_6379_out0;
wire v$RD_6380_out0;
wire v$RD_6381_out0;
wire v$RD_6382_out0;
wire v$RD_6383_out0;
wire v$RD_6384_out0;
wire v$RD_6385_out0;
wire v$RD_6386_out0;
wire v$RD_6387_out0;
wire v$RD_6388_out0;
wire v$RD_6389_out0;
wire v$RD_6390_out0;
wire v$RD_6391_out0;
wire v$RD_6392_out0;
wire v$RD_6393_out0;
wire v$RD_6394_out0;
wire v$RD_6395_out0;
wire v$RD_6396_out0;
wire v$RD_6397_out0;
wire v$RD_6398_out0;
wire v$RD_6399_out0;
wire v$RD_6400_out0;
wire v$RD_6401_out0;
wire v$RD_6402_out0;
wire v$RD_6403_out0;
wire v$RD_6404_out0;
wire v$RD_6405_out0;
wire v$RD_6406_out0;
wire v$RD_6407_out0;
wire v$RD_6408_out0;
wire v$RD_6409_out0;
wire v$RD_6410_out0;
wire v$RD_6411_out0;
wire v$RD_6412_out0;
wire v$RD_6413_out0;
wire v$RD_6414_out0;
wire v$RD_6415_out0;
wire v$RD_6416_out0;
wire v$RD_6417_out0;
wire v$RD_6418_out0;
wire v$RD_6419_out0;
wire v$RD_6420_out0;
wire v$RD_6421_out0;
wire v$RD_6422_out0;
wire v$RD_6423_out0;
wire v$RD_6424_out0;
wire v$RD_6425_out0;
wire v$RD_6426_out0;
wire v$RD_6427_out0;
wire v$RD_6428_out0;
wire v$RD_6429_out0;
wire v$RD_6430_out0;
wire v$RD_6431_out0;
wire v$RD_6432_out0;
wire v$RD_6433_out0;
wire v$RD_6434_out0;
wire v$RD_6435_out0;
wire v$RD_6436_out0;
wire v$RD_6437_out0;
wire v$RD_6438_out0;
wire v$RD_6439_out0;
wire v$RD_6440_out0;
wire v$RD_6441_out0;
wire v$RD_6442_out0;
wire v$RD_6443_out0;
wire v$RD_6444_out0;
wire v$RD_6445_out0;
wire v$RD_6446_out0;
wire v$RD_6447_out0;
wire v$RD_6448_out0;
wire v$RD_6449_out0;
wire v$RD_6450_out0;
wire v$RD_6451_out0;
wire v$RD_6452_out0;
wire v$RD_6453_out0;
wire v$RD_6454_out0;
wire v$RD_6455_out0;
wire v$RD_6456_out0;
wire v$RD_6457_out0;
wire v$RD_6458_out0;
wire v$RD_6459_out0;
wire v$RD_6460_out0;
wire v$RD_6461_out0;
wire v$RD_6462_out0;
wire v$RD_6463_out0;
wire v$RD_6464_out0;
wire v$RD_6465_out0;
wire v$RD_6466_out0;
wire v$RD_6467_out0;
wire v$RD_6468_out0;
wire v$RD_6469_out0;
wire v$RD_6470_out0;
wire v$RD_6471_out0;
wire v$RD_6472_out0;
wire v$RD_6473_out0;
wire v$RD_6474_out0;
wire v$RD_6475_out0;
wire v$RD_6476_out0;
wire v$RD_6477_out0;
wire v$RD_6478_out0;
wire v$RD_6479_out0;
wire v$RD_6480_out0;
wire v$RD_6481_out0;
wire v$RD_6482_out0;
wire v$RD_6483_out0;
wire v$RD_6484_out0;
wire v$RD_6485_out0;
wire v$RD_6486_out0;
wire v$RD_6487_out0;
wire v$RD_6488_out0;
wire v$RD_6489_out0;
wire v$RD_6490_out0;
wire v$RD_6491_out0;
wire v$RD_6492_out0;
wire v$RD_6493_out0;
wire v$RD_6494_out0;
wire v$RD_6495_out0;
wire v$RD_6496_out0;
wire v$RD_6497_out0;
wire v$RD_6498_out0;
wire v$RD_6499_out0;
wire v$RD_6500_out0;
wire v$RD_6501_out0;
wire v$RD_6502_out0;
wire v$RD_6503_out0;
wire v$RD_6504_out0;
wire v$RD_6505_out0;
wire v$RD_6506_out0;
wire v$RD_6507_out0;
wire v$RD_6508_out0;
wire v$RD_6509_out0;
wire v$RD_6510_out0;
wire v$RD_6511_out0;
wire v$RD_6512_out0;
wire v$RD_6513_out0;
wire v$RD_6514_out0;
wire v$RD_6515_out0;
wire v$RD_6516_out0;
wire v$RD_6517_out0;
wire v$RD_6518_out0;
wire v$RD_6519_out0;
wire v$RD_6520_out0;
wire v$RD_6521_out0;
wire v$RD_6522_out0;
wire v$RD_6523_out0;
wire v$RD_6524_out0;
wire v$RD_6525_out0;
wire v$RD_6526_out0;
wire v$RD_6527_out0;
wire v$RD_6528_out0;
wire v$RD_6529_out0;
wire v$RD_6530_out0;
wire v$RD_6531_out0;
wire v$RD_6532_out0;
wire v$RD_6533_out0;
wire v$RD_6534_out0;
wire v$RD_6535_out0;
wire v$RD_6536_out0;
wire v$RD_6537_out0;
wire v$RD_6538_out0;
wire v$RD_6539_out0;
wire v$RD_6540_out0;
wire v$RD_6541_out0;
wire v$RD_6542_out0;
wire v$RD_6543_out0;
wire v$RD_6544_out0;
wire v$RD_6545_out0;
wire v$RD_6546_out0;
wire v$RD_6547_out0;
wire v$RD_6548_out0;
wire v$RD_6549_out0;
wire v$RD_6550_out0;
wire v$RD_6551_out0;
wire v$RD_6552_out0;
wire v$RD_6553_out0;
wire v$RD_6554_out0;
wire v$RD_6555_out0;
wire v$RD_6556_out0;
wire v$RD_6557_out0;
wire v$RD_6558_out0;
wire v$RD_6559_out0;
wire v$RD_6560_out0;
wire v$RD_6561_out0;
wire v$RD_6562_out0;
wire v$RD_6563_out0;
wire v$RD_6564_out0;
wire v$RD_6565_out0;
wire v$RD_6566_out0;
wire v$RD_6567_out0;
wire v$RD_6568_out0;
wire v$RD_6569_out0;
wire v$RD_6570_out0;
wire v$RD_6571_out0;
wire v$RD_6572_out0;
wire v$RD_6573_out0;
wire v$RD_6574_out0;
wire v$RD_6575_out0;
wire v$RD_6576_out0;
wire v$RD_6577_out0;
wire v$RD_6578_out0;
wire v$RD_6579_out0;
wire v$RD_6580_out0;
wire v$RD_6581_out0;
wire v$RD_6582_out0;
wire v$RD_6583_out0;
wire v$RD_6584_out0;
wire v$RD_6585_out0;
wire v$RD_6586_out0;
wire v$RD_6587_out0;
wire v$RD_6588_out0;
wire v$RD_6589_out0;
wire v$RD_6590_out0;
wire v$RD_6591_out0;
wire v$RD_6592_out0;
wire v$RD_6593_out0;
wire v$RD_6594_out0;
wire v$RD_6595_out0;
wire v$RD_6596_out0;
wire v$RD_6597_out0;
wire v$RD_6598_out0;
wire v$RD_6599_out0;
wire v$RD_6600_out0;
wire v$RD_6601_out0;
wire v$RD_6602_out0;
wire v$RD_6603_out0;
wire v$RD_6604_out0;
wire v$RD_6605_out0;
wire v$RD_6606_out0;
wire v$RD_6607_out0;
wire v$RD_6608_out0;
wire v$RD_6609_out0;
wire v$RD_6610_out0;
wire v$RD_6611_out0;
wire v$RD_6612_out0;
wire v$RD_6613_out0;
wire v$RD_6614_out0;
wire v$RD_6615_out0;
wire v$RD_6616_out0;
wire v$RD_6617_out0;
wire v$RD_6618_out0;
wire v$RD_6619_out0;
wire v$RD_6620_out0;
wire v$RD_6621_out0;
wire v$RD_6622_out0;
wire v$RD_6623_out0;
wire v$RD_6624_out0;
wire v$RD_6625_out0;
wire v$RD_6626_out0;
wire v$RD_6627_out0;
wire v$RD_6628_out0;
wire v$RD_6629_out0;
wire v$RD_6630_out0;
wire v$RD_6631_out0;
wire v$RD_6632_out0;
wire v$RD_6633_out0;
wire v$RD_6634_out0;
wire v$RD_6635_out0;
wire v$RD_6636_out0;
wire v$RD_6637_out0;
wire v$RD_6638_out0;
wire v$RD_6639_out0;
wire v$RD_6640_out0;
wire v$RD_6641_out0;
wire v$RD_6642_out0;
wire v$RD_6643_out0;
wire v$RD_6644_out0;
wire v$RD_6645_out0;
wire v$RD_6646_out0;
wire v$RD_6647_out0;
wire v$RD_6648_out0;
wire v$RD_6649_out0;
wire v$RD_6650_out0;
wire v$RD_6651_out0;
wire v$RD_6652_out0;
wire v$RD_6653_out0;
wire v$RD_6654_out0;
wire v$RD_6655_out0;
wire v$RD_6656_out0;
wire v$RD_6657_out0;
wire v$RD_6658_out0;
wire v$RD_6659_out0;
wire v$RD_6660_out0;
wire v$RD_6661_out0;
wire v$RD_6662_out0;
wire v$RD_6663_out0;
wire v$RD_6664_out0;
wire v$RD_6665_out0;
wire v$RD_6666_out0;
wire v$RD_6667_out0;
wire v$RD_6668_out0;
wire v$RD_6669_out0;
wire v$RD_6670_out0;
wire v$RD_6671_out0;
wire v$RD_6672_out0;
wire v$RD_6673_out0;
wire v$RD_6674_out0;
wire v$RD_6675_out0;
wire v$RD_6676_out0;
wire v$RD_6677_out0;
wire v$RD_6678_out0;
wire v$RD_6679_out0;
wire v$RD_6680_out0;
wire v$RD_6681_out0;
wire v$RD_6682_out0;
wire v$RD_6683_out0;
wire v$RD_6684_out0;
wire v$RD_6685_out0;
wire v$RD_6686_out0;
wire v$RD_6687_out0;
wire v$RD_6688_out0;
wire v$RD_6689_out0;
wire v$RD_6690_out0;
wire v$RD_6691_out0;
wire v$RD_6692_out0;
wire v$RD_6693_out0;
wire v$RD_6694_out0;
wire v$RD_6695_out0;
wire v$RD_6696_out0;
wire v$RD_6697_out0;
wire v$RD_6698_out0;
wire v$RD_6699_out0;
wire v$RD_6700_out0;
wire v$RD_6701_out0;
wire v$RD_6702_out0;
wire v$RD_6703_out0;
wire v$RD_6704_out0;
wire v$RD_6705_out0;
wire v$RD_6706_out0;
wire v$RD_6707_out0;
wire v$RD_6708_out0;
wire v$RD_6709_out0;
wire v$RD_6710_out0;
wire v$RD_6711_out0;
wire v$RD_6712_out0;
wire v$RD_6713_out0;
wire v$RD_6714_out0;
wire v$RD_6715_out0;
wire v$RD_6716_out0;
wire v$RD_6717_out0;
wire v$RD_6718_out0;
wire v$RD_6719_out0;
wire v$RD_6720_out0;
wire v$RD_6721_out0;
wire v$RD_6722_out0;
wire v$RD_6723_out0;
wire v$RD_6724_out0;
wire v$RD_6725_out0;
wire v$RD_6726_out0;
wire v$RD_6727_out0;
wire v$RD_6728_out0;
wire v$RD_6729_out0;
wire v$RD_6730_out0;
wire v$RD_6731_out0;
wire v$RD_6732_out0;
wire v$RD_6733_out0;
wire v$RD_6734_out0;
wire v$RD_6735_out0;
wire v$RD_6736_out0;
wire v$RD_6737_out0;
wire v$RD_6738_out0;
wire v$RD_6739_out0;
wire v$RD_6740_out0;
wire v$RD_6741_out0;
wire v$RD_6742_out0;
wire v$RD_6743_out0;
wire v$RD_6744_out0;
wire v$RD_6745_out0;
wire v$RD_6746_out0;
wire v$RD_6747_out0;
wire v$RD_6748_out0;
wire v$RD_6749_out0;
wire v$RD_6750_out0;
wire v$RD_6751_out0;
wire v$RD_6752_out0;
wire v$RD_6753_out0;
wire v$RD_6754_out0;
wire v$RD_6755_out0;
wire v$RD_6756_out0;
wire v$RD_6757_out0;
wire v$RD_6758_out0;
wire v$RD_6759_out0;
wire v$RD_6760_out0;
wire v$RD_6761_out0;
wire v$RD_6762_out0;
wire v$RD_6763_out0;
wire v$RD_6764_out0;
wire v$RD_6765_out0;
wire v$RD_6766_out0;
wire v$RD_6767_out0;
wire v$RD_6768_out0;
wire v$RD_6769_out0;
wire v$RD_6770_out0;
wire v$RD_6771_out0;
wire v$RD_6772_out0;
wire v$RD_6773_out0;
wire v$RD_6774_out0;
wire v$RD_6775_out0;
wire v$RD_6776_out0;
wire v$RD_6777_out0;
wire v$RD_6778_out0;
wire v$RD_6779_out0;
wire v$RD_6780_out0;
wire v$RD_6781_out0;
wire v$RD_6782_out0;
wire v$RD_6783_out0;
wire v$RD_6784_out0;
wire v$RD_6785_out0;
wire v$RD_6786_out0;
wire v$RD_6787_out0;
wire v$RD_6788_out0;
wire v$RD_6789_out0;
wire v$RD_7187_out0;
wire v$RD_7188_out0;
wire v$RD_7189_out0;
wire v$RD_7190_out0;
wire v$RD_7191_out0;
wire v$RD_7192_out0;
wire v$RD_7193_out0;
wire v$RD_7194_out0;
wire v$RD_7195_out0;
wire v$RD_7196_out0;
wire v$RD_7197_out0;
wire v$RD_7198_out0;
wire v$RD_7199_out0;
wire v$RD_7200_out0;
wire v$RD_7201_out0;
wire v$RD_7202_out0;
wire v$RD_7203_out0;
wire v$RD_7204_out0;
wire v$RD_7205_out0;
wire v$RD_7206_out0;
wire v$RD_7207_out0;
wire v$RD_7208_out0;
wire v$RD_7209_out0;
wire v$RD_7210_out0;
wire v$RD_7211_out0;
wire v$RD_7212_out0;
wire v$RD_7213_out0;
wire v$RD_7214_out0;
wire v$RD_7215_out0;
wire v$RD_7216_out0;
wire v$RD_7217_out0;
wire v$RD_7218_out0;
wire v$RD_7219_out0;
wire v$RD_7220_out0;
wire v$RD_7221_out0;
wire v$RD_7222_out0;
wire v$RD_7223_out0;
wire v$RD_7224_out0;
wire v$RD_7225_out0;
wire v$RD_7226_out0;
wire v$RD_7227_out0;
wire v$RD_7228_out0;
wire v$RD_7229_out0;
wire v$RD_7230_out0;
wire v$RD_7231_out0;
wire v$RD_7232_out0;
wire v$RD_7233_out0;
wire v$RD_7234_out0;
wire v$RD_7235_out0;
wire v$RD_7236_out0;
wire v$RD_7237_out0;
wire v$RD_7238_out0;
wire v$RD_7239_out0;
wire v$RD_7240_out0;
wire v$RD_7241_out0;
wire v$RD_7242_out0;
wire v$RD_7243_out0;
wire v$RD_7244_out0;
wire v$RD_7245_out0;
wire v$RD_7246_out0;
wire v$RD_7247_out0;
wire v$RD_7248_out0;
wire v$RD_7249_out0;
wire v$RD_7250_out0;
wire v$RD_7251_out0;
wire v$RD_7252_out0;
wire v$RD_7253_out0;
wire v$RD_7254_out0;
wire v$RD_7255_out0;
wire v$RD_7256_out0;
wire v$RD_7257_out0;
wire v$RD_7258_out0;
wire v$RD_7259_out0;
wire v$RD_7260_out0;
wire v$RD_7261_out0;
wire v$RD_7262_out0;
wire v$RD_7263_out0;
wire v$RD_7264_out0;
wire v$RD_7265_out0;
wire v$RD_7266_out0;
wire v$RD_7267_out0;
wire v$RD_7268_out0;
wire v$RD_7269_out0;
wire v$RD_7270_out0;
wire v$RD_7271_out0;
wire v$RD_7272_out0;
wire v$RD_7273_out0;
wire v$RD_7274_out0;
wire v$RD_7275_out0;
wire v$RD_7276_out0;
wire v$RD_7277_out0;
wire v$RD_7278_out0;
wire v$RD_7279_out0;
wire v$RD_7280_out0;
wire v$RD_7281_out0;
wire v$RD_7282_out0;
wire v$RD_7283_out0;
wire v$RD_7284_out0;
wire v$RD_7285_out0;
wire v$RD_7286_out0;
wire v$RD_7287_out0;
wire v$RD_7288_out0;
wire v$RD_7289_out0;
wire v$RD_7290_out0;
wire v$RD_7291_out0;
wire v$RD_7292_out0;
wire v$RD_7293_out0;
wire v$RD_7294_out0;
wire v$RD_7295_out0;
wire v$RD_7296_out0;
wire v$RD_7297_out0;
wire v$RD_7298_out0;
wire v$RD_7299_out0;
wire v$RD_7300_out0;
wire v$RD_7301_out0;
wire v$RD_7302_out0;
wire v$RD_7303_out0;
wire v$RD_7304_out0;
wire v$RD_7305_out0;
wire v$RD_7306_out0;
wire v$RD_7307_out0;
wire v$RD_7308_out0;
wire v$RD_7309_out0;
wire v$RD_7310_out0;
wire v$RD_7311_out0;
wire v$RD_7312_out0;
wire v$RD_7313_out0;
wire v$RD_7314_out0;
wire v$RD_7315_out0;
wire v$RD_7316_out0;
wire v$RD_7317_out0;
wire v$RD_7318_out0;
wire v$RD_7319_out0;
wire v$RD_7320_out0;
wire v$RD_7321_out0;
wire v$RD_7322_out0;
wire v$RD_7323_out0;
wire v$RD_7324_out0;
wire v$RD_7325_out0;
wire v$RD_7326_out0;
wire v$RD_7327_out0;
wire v$RD_7328_out0;
wire v$RD_7329_out0;
wire v$RD_7330_out0;
wire v$RD_7331_out0;
wire v$RD_7332_out0;
wire v$RD_7333_out0;
wire v$RD_7334_out0;
wire v$RD_7335_out0;
wire v$RD_7336_out0;
wire v$RD_7337_out0;
wire v$RD_7338_out0;
wire v$RD_7339_out0;
wire v$RD_7340_out0;
wire v$RD_7341_out0;
wire v$RD_7342_out0;
wire v$RD_7343_out0;
wire v$RD_7344_out0;
wire v$RD_7345_out0;
wire v$RD_7346_out0;
wire v$RD_7347_out0;
wire v$RD_7348_out0;
wire v$RD_7349_out0;
wire v$RD_7350_out0;
wire v$RD_7351_out0;
wire v$RD_7352_out0;
wire v$RD_7353_out0;
wire v$RD_7354_out0;
wire v$RD_7355_out0;
wire v$RD_7356_out0;
wire v$RD_7357_out0;
wire v$RD_7358_out0;
wire v$RD_7359_out0;
wire v$RD_7360_out0;
wire v$RD_7361_out0;
wire v$RD_7362_out0;
wire v$RD_7363_out0;
wire v$RD_7364_out0;
wire v$RD_7365_out0;
wire v$RD_7366_out0;
wire v$RD_7367_out0;
wire v$RD_7368_out0;
wire v$RD_7369_out0;
wire v$RD_7370_out0;
wire v$RD_7371_out0;
wire v$RD_7372_out0;
wire v$RD_7373_out0;
wire v$RD_7374_out0;
wire v$RD_7375_out0;
wire v$RD_7376_out0;
wire v$RD_7377_out0;
wire v$RD_7378_out0;
wire v$RD_7379_out0;
wire v$RD_7380_out0;
wire v$RD_7381_out0;
wire v$RD_7382_out0;
wire v$RD_7383_out0;
wire v$RD_7384_out0;
wire v$RD_7385_out0;
wire v$RD_7386_out0;
wire v$RD_7387_out0;
wire v$RD_7388_out0;
wire v$RD_7389_out0;
wire v$RD_7390_out0;
wire v$RD_7391_out0;
wire v$RD_7392_out0;
wire v$RD_7393_out0;
wire v$RD_7394_out0;
wire v$RD_7395_out0;
wire v$RD_7396_out0;
wire v$RD_7397_out0;
wire v$RD_7398_out0;
wire v$RD_7399_out0;
wire v$RD_7400_out0;
wire v$RD_7401_out0;
wire v$RD_7402_out0;
wire v$RD_7403_out0;
wire v$RD_7404_out0;
wire v$RD_7405_out0;
wire v$RD_7406_out0;
wire v$RD_7407_out0;
wire v$RD_7408_out0;
wire v$RD_7409_out0;
wire v$RD_7410_out0;
wire v$RD_7411_out0;
wire v$RD_7412_out0;
wire v$RD_7413_out0;
wire v$RD_7414_out0;
wire v$RD_7415_out0;
wire v$RD_7416_out0;
wire v$RD_7417_out0;
wire v$RD_7418_out0;
wire v$RD_7419_out0;
wire v$RD_7420_out0;
wire v$RD_7421_out0;
wire v$RD_7422_out0;
wire v$RD_7423_out0;
wire v$RD_7424_out0;
wire v$RD_7425_out0;
wire v$RD_7426_out0;
wire v$RD_7427_out0;
wire v$RD_7428_out0;
wire v$RD_7429_out0;
wire v$RD_7430_out0;
wire v$RD_7431_out0;
wire v$RD_7432_out0;
wire v$RD_7433_out0;
wire v$RD_7434_out0;
wire v$RD_7435_out0;
wire v$RD_7436_out0;
wire v$RD_7437_out0;
wire v$RD_7438_out0;
wire v$RD_7439_out0;
wire v$RD_7440_out0;
wire v$RD_7441_out0;
wire v$RD_7442_out0;
wire v$RD_7443_out0;
wire v$RD_7444_out0;
wire v$RD_7445_out0;
wire v$RD_7446_out0;
wire v$RD_7447_out0;
wire v$RD_7448_out0;
wire v$RD_7449_out0;
wire v$RD_7450_out0;
wire v$RD_7451_out0;
wire v$RD_7452_out0;
wire v$RD_7453_out0;
wire v$RD_7454_out0;
wire v$RD_7455_out0;
wire v$RD_7456_out0;
wire v$RD_7457_out0;
wire v$RD_7458_out0;
wire v$RD_7459_out0;
wire v$RD_7460_out0;
wire v$RD_7461_out0;
wire v$RD_7462_out0;
wire v$RD_7463_out0;
wire v$RD_7464_out0;
wire v$RD_7465_out0;
wire v$RD_7466_out0;
wire v$RD_7467_out0;
wire v$RD_7468_out0;
wire v$RD_7469_out0;
wire v$RD_7470_out0;
wire v$RD_7471_out0;
wire v$RD_7472_out0;
wire v$RD_7473_out0;
wire v$RD_7474_out0;
wire v$RD_7475_out0;
wire v$RD_7476_out0;
wire v$RD_7477_out0;
wire v$RD_7478_out0;
wire v$RD_7479_out0;
wire v$RD_7480_out0;
wire v$RD_7481_out0;
wire v$RD_7482_out0;
wire v$RD_7483_out0;
wire v$RD_7484_out0;
wire v$RD_7485_out0;
wire v$RD_7486_out0;
wire v$RD_7487_out0;
wire v$RD_7488_out0;
wire v$RD_7489_out0;
wire v$RD_7490_out0;
wire v$RD_7491_out0;
wire v$RD_7492_out0;
wire v$RD_7493_out0;
wire v$RD_7494_out0;
wire v$RD_7495_out0;
wire v$RD_7496_out0;
wire v$RD_7497_out0;
wire v$RD_7498_out0;
wire v$RD_7499_out0;
wire v$RD_7500_out0;
wire v$RD_7501_out0;
wire v$RD_7502_out0;
wire v$RD_7503_out0;
wire v$RD_7504_out0;
wire v$RD_7505_out0;
wire v$RD_7506_out0;
wire v$RD_7507_out0;
wire v$RD_7508_out0;
wire v$RD_7509_out0;
wire v$RD_7510_out0;
wire v$RD_7511_out0;
wire v$RD_7512_out0;
wire v$RD_7513_out0;
wire v$RD_7514_out0;
wire v$RD_7515_out0;
wire v$RD_7516_out0;
wire v$RD_7517_out0;
wire v$RD_7518_out0;
wire v$RD_7519_out0;
wire v$RD_7520_out0;
wire v$RD_7521_out0;
wire v$RD_7522_out0;
wire v$RD_7523_out0;
wire v$RD_7524_out0;
wire v$RD_7525_out0;
wire v$RD_7526_out0;
wire v$RD_7527_out0;
wire v$RD_7528_out0;
wire v$RD_7529_out0;
wire v$RD_7530_out0;
wire v$RD_7531_out0;
wire v$RD_7532_out0;
wire v$RD_7533_out0;
wire v$RD_7534_out0;
wire v$RD_7535_out0;
wire v$RD_7536_out0;
wire v$RD_7537_out0;
wire v$RD_7538_out0;
wire v$RD_7539_out0;
wire v$RD_7540_out0;
wire v$RD_7541_out0;
wire v$RD_7542_out0;
wire v$RD_7543_out0;
wire v$RD_7544_out0;
wire v$RD_7545_out0;
wire v$RD_7546_out0;
wire v$RD_7547_out0;
wire v$RD_7548_out0;
wire v$RD_7549_out0;
wire v$RD_7550_out0;
wire v$RD_7551_out0;
wire v$RD_7552_out0;
wire v$RD_7553_out0;
wire v$RD_7554_out0;
wire v$RD_7555_out0;
wire v$RD_7556_out0;
wire v$RD_7557_out0;
wire v$RD_7558_out0;
wire v$RD_7559_out0;
wire v$RD_7560_out0;
wire v$RD_7561_out0;
wire v$RD_7562_out0;
wire v$RD_7563_out0;
wire v$RD_7564_out0;
wire v$RD_7565_out0;
wire v$RD_7566_out0;
wire v$RD_7567_out0;
wire v$RD_7568_out0;
wire v$RD_7569_out0;
wire v$RD_7570_out0;
wire v$RD_7571_out0;
wire v$RD_7572_out0;
wire v$RD_7573_out0;
wire v$RD_7574_out0;
wire v$RD_7575_out0;
wire v$RD_7576_out0;
wire v$RD_7577_out0;
wire v$RD_7578_out0;
wire v$RD_7579_out0;
wire v$RD_7580_out0;
wire v$RD_7581_out0;
wire v$RD_7582_out0;
wire v$RD_7583_out0;
wire v$RD_7584_out0;
wire v$RD_7585_out0;
wire v$RD_7586_out0;
wire v$RD_7587_out0;
wire v$RD_7588_out0;
wire v$RD_7589_out0;
wire v$RD_7590_out0;
wire v$RD_7591_out0;
wire v$RD_7592_out0;
wire v$RD_7593_out0;
wire v$RD_7594_out0;
wire v$RD_7595_out0;
wire v$RD_7596_out0;
wire v$RD_7597_out0;
wire v$RD_7598_out0;
wire v$RD_7599_out0;
wire v$RD_7600_out0;
wire v$RD_7601_out0;
wire v$RD_7602_out0;
wire v$RD_7603_out0;
wire v$RD_7604_out0;
wire v$RD_7605_out0;
wire v$RD_7606_out0;
wire v$RD_7607_out0;
wire v$RD_7608_out0;
wire v$RD_7609_out0;
wire v$RD_7610_out0;
wire v$RD_7611_out0;
wire v$RD_7612_out0;
wire v$RD_7613_out0;
wire v$RD_7614_out0;
wire v$RD_7615_out0;
wire v$RD_7616_out0;
wire v$RD_7617_out0;
wire v$RD_7618_out0;
wire v$RD_7619_out0;
wire v$RD_7620_out0;
wire v$RD_7621_out0;
wire v$RD_7622_out0;
wire v$RD_7623_out0;
wire v$RD_7624_out0;
wire v$RD_7625_out0;
wire v$RD_7626_out0;
wire v$RD_7627_out0;
wire v$RD_7628_out0;
wire v$RD_7629_out0;
wire v$RD_7630_out0;
wire v$RD_7631_out0;
wire v$RD_7632_out0;
wire v$RD_7633_out0;
wire v$RD_7634_out0;
wire v$REN0_11136_out0;
wire v$REN1_6874_out0;
wire v$RESET_11174_out0;
wire v$RESET_11175_out0;
wire v$RESET_11176_out0;
wire v$RESET_11177_out0;
wire v$RESET_11178_out0;
wire v$RESET_11179_out0;
wire v$RESET_11180_out0;
wire v$RESET_11181_out0;
wire v$RESET_11182_out0;
wire v$RESET_11183_out0;
wire v$RESET_11184_out0;
wire v$RESET_11185_out0;
wire v$RESET_11186_out0;
wire v$RESET_11187_out0;
wire v$RESET_11188_out0;
wire v$RESET_11189_out0;
wire v$RM_11302_out0;
wire v$RM_11303_out0;
wire v$RM_11304_out0;
wire v$RM_11305_out0;
wire v$RM_11306_out0;
wire v$RM_11307_out0;
wire v$RM_11308_out0;
wire v$RM_11309_out0;
wire v$RM_11310_out0;
wire v$RM_11311_out0;
wire v$RM_11312_out0;
wire v$RM_11313_out0;
wire v$RM_11314_out0;
wire v$RM_11315_out0;
wire v$RM_11316_out0;
wire v$RM_11317_out0;
wire v$RM_11318_out0;
wire v$RM_11319_out0;
wire v$RM_11320_out0;
wire v$RM_11321_out0;
wire v$RM_11322_out0;
wire v$RM_11323_out0;
wire v$RM_11324_out0;
wire v$RM_11325_out0;
wire v$RM_11326_out0;
wire v$RM_11327_out0;
wire v$RM_11328_out0;
wire v$RM_11329_out0;
wire v$RM_11330_out0;
wire v$RM_11331_out0;
wire v$RM_11332_out0;
wire v$RM_11333_out0;
wire v$RM_11334_out0;
wire v$RM_11335_out0;
wire v$RM_11336_out0;
wire v$RM_11337_out0;
wire v$RM_11338_out0;
wire v$RM_11339_out0;
wire v$RM_11340_out0;
wire v$RM_11341_out0;
wire v$RM_11342_out0;
wire v$RM_11343_out0;
wire v$RM_11344_out0;
wire v$RM_11345_out0;
wire v$RM_11346_out0;
wire v$RM_11347_out0;
wire v$RM_11348_out0;
wire v$RM_11349_out0;
wire v$RM_11350_out0;
wire v$RM_11351_out0;
wire v$RM_11352_out0;
wire v$RM_11353_out0;
wire v$RM_11354_out0;
wire v$RM_11355_out0;
wire v$RM_11356_out0;
wire v$RM_11357_out0;
wire v$RM_11358_out0;
wire v$RM_11359_out0;
wire v$RM_11360_out0;
wire v$RM_11361_out0;
wire v$RM_11362_out0;
wire v$RM_11363_out0;
wire v$RM_11364_out0;
wire v$RM_11365_out0;
wire v$RM_11366_out0;
wire v$RM_11367_out0;
wire v$RM_11368_out0;
wire v$RM_11369_out0;
wire v$RM_11370_out0;
wire v$RM_11371_out0;
wire v$RM_11372_out0;
wire v$RM_11373_out0;
wire v$RM_11374_out0;
wire v$RM_11375_out0;
wire v$RM_11376_out0;
wire v$RM_11377_out0;
wire v$RM_11378_out0;
wire v$RM_11379_out0;
wire v$RM_11380_out0;
wire v$RM_11381_out0;
wire v$RM_11382_out0;
wire v$RM_11383_out0;
wire v$RM_11384_out0;
wire v$RM_11385_out0;
wire v$RM_11386_out0;
wire v$RM_11387_out0;
wire v$RM_11388_out0;
wire v$RM_11389_out0;
wire v$RM_11390_out0;
wire v$RM_11391_out0;
wire v$RM_11392_out0;
wire v$RM_11393_out0;
wire v$RM_11394_out0;
wire v$RM_11395_out0;
wire v$RM_11396_out0;
wire v$RM_11397_out0;
wire v$RM_11398_out0;
wire v$RM_11399_out0;
wire v$RM_11400_out0;
wire v$RM_11401_out0;
wire v$RM_11402_out0;
wire v$RM_11403_out0;
wire v$RM_11404_out0;
wire v$RM_11405_out0;
wire v$RM_11406_out0;
wire v$RM_11407_out0;
wire v$RM_11408_out0;
wire v$RM_11409_out0;
wire v$RM_11410_out0;
wire v$RM_11411_out0;
wire v$RM_11412_out0;
wire v$RM_11413_out0;
wire v$RM_11414_out0;
wire v$RM_11415_out0;
wire v$RM_11416_out0;
wire v$RM_11417_out0;
wire v$RM_11418_out0;
wire v$RM_11419_out0;
wire v$RM_11420_out0;
wire v$RM_11421_out0;
wire v$RM_11422_out0;
wire v$RM_11423_out0;
wire v$RM_11424_out0;
wire v$RM_11425_out0;
wire v$RM_11426_out0;
wire v$RM_11427_out0;
wire v$RM_11428_out0;
wire v$RM_11429_out0;
wire v$RM_11430_out0;
wire v$RM_11431_out0;
wire v$RM_11432_out0;
wire v$RM_11433_out0;
wire v$RM_11434_out0;
wire v$RM_11435_out0;
wire v$RM_11436_out0;
wire v$RM_11437_out0;
wire v$RM_11438_out0;
wire v$RM_11439_out0;
wire v$RM_11440_out0;
wire v$RM_11441_out0;
wire v$RM_11442_out0;
wire v$RM_11443_out0;
wire v$RM_11444_out0;
wire v$RM_11445_out0;
wire v$RM_11446_out0;
wire v$RM_11447_out0;
wire v$RM_11448_out0;
wire v$RM_11449_out0;
wire v$RM_11450_out0;
wire v$RM_11451_out0;
wire v$RM_11452_out0;
wire v$RM_11453_out0;
wire v$RM_11454_out0;
wire v$RM_11455_out0;
wire v$RM_11456_out0;
wire v$RM_11457_out0;
wire v$RM_11458_out0;
wire v$RM_11459_out0;
wire v$RM_11460_out0;
wire v$RM_11461_out0;
wire v$RM_11462_out0;
wire v$RM_11463_out0;
wire v$RM_11464_out0;
wire v$RM_11465_out0;
wire v$RM_11466_out0;
wire v$RM_11467_out0;
wire v$RM_11468_out0;
wire v$RM_11469_out0;
wire v$RM_11470_out0;
wire v$RM_11471_out0;
wire v$RM_11472_out0;
wire v$RM_11473_out0;
wire v$RM_11474_out0;
wire v$RM_11475_out0;
wire v$RM_11476_out0;
wire v$RM_11477_out0;
wire v$RM_11478_out0;
wire v$RM_11479_out0;
wire v$RM_11480_out0;
wire v$RM_11481_out0;
wire v$RM_11482_out0;
wire v$RM_11483_out0;
wire v$RM_11484_out0;
wire v$RM_11485_out0;
wire v$RM_11486_out0;
wire v$RM_11487_out0;
wire v$RM_11488_out0;
wire v$RM_11489_out0;
wire v$RM_11490_out0;
wire v$RM_11491_out0;
wire v$RM_11492_out0;
wire v$RM_11493_out0;
wire v$RM_11494_out0;
wire v$RM_11495_out0;
wire v$RM_11496_out0;
wire v$RM_11497_out0;
wire v$RM_11498_out0;
wire v$RM_11499_out0;
wire v$RM_11500_out0;
wire v$RM_11501_out0;
wire v$RM_11502_out0;
wire v$RM_11503_out0;
wire v$RM_11504_out0;
wire v$RM_11505_out0;
wire v$RM_11506_out0;
wire v$RM_11507_out0;
wire v$RM_11508_out0;
wire v$RM_11509_out0;
wire v$RM_11510_out0;
wire v$RM_11511_out0;
wire v$RM_11512_out0;
wire v$RM_11513_out0;
wire v$RM_11514_out0;
wire v$RM_11515_out0;
wire v$RM_11516_out0;
wire v$RM_11517_out0;
wire v$RM_11518_out0;
wire v$RM_11519_out0;
wire v$RM_11520_out0;
wire v$RM_11521_out0;
wire v$RM_11522_out0;
wire v$RM_11523_out0;
wire v$RM_11524_out0;
wire v$RM_11525_out0;
wire v$RM_11526_out0;
wire v$RM_11527_out0;
wire v$RM_11528_out0;
wire v$RM_11529_out0;
wire v$RM_11530_out0;
wire v$RM_11531_out0;
wire v$RM_11532_out0;
wire v$RM_11533_out0;
wire v$RM_11534_out0;
wire v$RM_11535_out0;
wire v$RM_11536_out0;
wire v$RM_11537_out0;
wire v$RM_11538_out0;
wire v$RM_11539_out0;
wire v$RM_11540_out0;
wire v$RM_11541_out0;
wire v$RM_11542_out0;
wire v$RM_11543_out0;
wire v$RM_11544_out0;
wire v$RM_11545_out0;
wire v$RM_11546_out0;
wire v$RM_11547_out0;
wire v$RM_11548_out0;
wire v$RM_11549_out0;
wire v$RM_11550_out0;
wire v$RM_11551_out0;
wire v$RM_11552_out0;
wire v$RM_11553_out0;
wire v$RM_11554_out0;
wire v$RM_11555_out0;
wire v$RM_11556_out0;
wire v$RM_11557_out0;
wire v$RM_11558_out0;
wire v$RM_11559_out0;
wire v$RM_11560_out0;
wire v$RM_11561_out0;
wire v$RM_11562_out0;
wire v$RM_11563_out0;
wire v$RM_11564_out0;
wire v$RM_11565_out0;
wire v$RM_11566_out0;
wire v$RM_11567_out0;
wire v$RM_11568_out0;
wire v$RM_11569_out0;
wire v$RM_11570_out0;
wire v$RM_11571_out0;
wire v$RM_11572_out0;
wire v$RM_11573_out0;
wire v$RM_11574_out0;
wire v$RM_11575_out0;
wire v$RM_11576_out0;
wire v$RM_11577_out0;
wire v$RM_11578_out0;
wire v$RM_11579_out0;
wire v$RM_11580_out0;
wire v$RM_11581_out0;
wire v$RM_11582_out0;
wire v$RM_11583_out0;
wire v$RM_11584_out0;
wire v$RM_11585_out0;
wire v$RM_11586_out0;
wire v$RM_11587_out0;
wire v$RM_11588_out0;
wire v$RM_11589_out0;
wire v$RM_11590_out0;
wire v$RM_11591_out0;
wire v$RM_11592_out0;
wire v$RM_11593_out0;
wire v$RM_11594_out0;
wire v$RM_11595_out0;
wire v$RM_11596_out0;
wire v$RM_11597_out0;
wire v$RM_11598_out0;
wire v$RM_11599_out0;
wire v$RM_11600_out0;
wire v$RM_11601_out0;
wire v$RM_11602_out0;
wire v$RM_11603_out0;
wire v$RM_11604_out0;
wire v$RM_11605_out0;
wire v$RM_11606_out0;
wire v$RM_11607_out0;
wire v$RM_11608_out0;
wire v$RM_11609_out0;
wire v$RM_11610_out0;
wire v$RM_11611_out0;
wire v$RM_11612_out0;
wire v$RM_11613_out0;
wire v$RM_11614_out0;
wire v$RM_11615_out0;
wire v$RM_11616_out0;
wire v$RM_11617_out0;
wire v$RM_11618_out0;
wire v$RM_11619_out0;
wire v$RM_11620_out0;
wire v$RM_11621_out0;
wire v$RM_11622_out0;
wire v$RM_11623_out0;
wire v$RM_11624_out0;
wire v$RM_11625_out0;
wire v$RM_11626_out0;
wire v$RM_11627_out0;
wire v$RM_11628_out0;
wire v$RM_11629_out0;
wire v$RM_11630_out0;
wire v$RM_11631_out0;
wire v$RM_11632_out0;
wire v$RM_11633_out0;
wire v$RM_11634_out0;
wire v$RM_11635_out0;
wire v$RM_11636_out0;
wire v$RM_11637_out0;
wire v$RM_11638_out0;
wire v$RM_11639_out0;
wire v$RM_11640_out0;
wire v$RM_11641_out0;
wire v$RM_11642_out0;
wire v$RM_11643_out0;
wire v$RM_11644_out0;
wire v$RM_11645_out0;
wire v$RM_11646_out0;
wire v$RM_11647_out0;
wire v$RM_11648_out0;
wire v$RM_11649_out0;
wire v$RM_11650_out0;
wire v$RM_11651_out0;
wire v$RM_11652_out0;
wire v$RM_11653_out0;
wire v$RM_11654_out0;
wire v$RM_11655_out0;
wire v$RM_11656_out0;
wire v$RM_11657_out0;
wire v$RM_11658_out0;
wire v$RM_11659_out0;
wire v$RM_11660_out0;
wire v$RM_11661_out0;
wire v$RM_11662_out0;
wire v$RM_11663_out0;
wire v$RM_11664_out0;
wire v$RM_11665_out0;
wire v$RM_11666_out0;
wire v$RM_11667_out0;
wire v$RM_11668_out0;
wire v$RM_11669_out0;
wire v$RM_11670_out0;
wire v$RM_11671_out0;
wire v$RM_11672_out0;
wire v$RM_11673_out0;
wire v$RM_11674_out0;
wire v$RM_11675_out0;
wire v$RM_11676_out0;
wire v$RM_11677_out0;
wire v$RM_11678_out0;
wire v$RM_11679_out0;
wire v$RM_11680_out0;
wire v$RM_11681_out0;
wire v$RM_11682_out0;
wire v$RM_11683_out0;
wire v$RM_11684_out0;
wire v$RM_11685_out0;
wire v$RM_11686_out0;
wire v$RM_11687_out0;
wire v$RM_11688_out0;
wire v$RM_11689_out0;
wire v$RM_11690_out0;
wire v$RM_11691_out0;
wire v$RM_11692_out0;
wire v$RM_11693_out0;
wire v$RM_11694_out0;
wire v$RM_11695_out0;
wire v$RM_11696_out0;
wire v$RM_11697_out0;
wire v$RM_11698_out0;
wire v$RM_11699_out0;
wire v$RM_11700_out0;
wire v$RM_11701_out0;
wire v$RM_11702_out0;
wire v$RM_11703_out0;
wire v$RM_11704_out0;
wire v$RM_11705_out0;
wire v$RM_11706_out0;
wire v$RM_11707_out0;
wire v$RM_11708_out0;
wire v$RM_11709_out0;
wire v$RM_11710_out0;
wire v$RM_11711_out0;
wire v$RM_11712_out0;
wire v$RM_11713_out0;
wire v$RM_11714_out0;
wire v$RM_11715_out0;
wire v$RM_11716_out0;
wire v$RM_11717_out0;
wire v$RM_11718_out0;
wire v$RM_11719_out0;
wire v$RM_11720_out0;
wire v$RM_11721_out0;
wire v$RM_11722_out0;
wire v$RM_11723_out0;
wire v$RM_11724_out0;
wire v$RM_11725_out0;
wire v$RM_11726_out0;
wire v$RM_11727_out0;
wire v$RM_11728_out0;
wire v$RM_11729_out0;
wire v$RM_11730_out0;
wire v$RM_11731_out0;
wire v$RM_11732_out0;
wire v$RM_11733_out0;
wire v$RM_11734_out0;
wire v$RM_11735_out0;
wire v$RM_11736_out0;
wire v$RM_11737_out0;
wire v$RM_11738_out0;
wire v$RM_11739_out0;
wire v$RM_11740_out0;
wire v$RM_11741_out0;
wire v$RM_11742_out0;
wire v$RM_11743_out0;
wire v$RM_11744_out0;
wire v$RM_11745_out0;
wire v$RM_11746_out0;
wire v$RM_11747_out0;
wire v$RM_11748_out0;
wire v$RM_11749_out0;
wire v$RM_11750_out0;
wire v$RM_11751_out0;
wire v$RM_11752_out0;
wire v$RM_11753_out0;
wire v$RM_11754_out0;
wire v$RM_11755_out0;
wire v$RM_11756_out0;
wire v$RM_11757_out0;
wire v$RM_11758_out0;
wire v$RM_11759_out0;
wire v$RM_11760_out0;
wire v$RM_11761_out0;
wire v$RM_11762_out0;
wire v$RM_11763_out0;
wire v$RM_11764_out0;
wire v$RM_11765_out0;
wire v$RM_11766_out0;
wire v$RM_11767_out0;
wire v$RM_11768_out0;
wire v$RM_11769_out0;
wire v$RM_11770_out0;
wire v$RM_11771_out0;
wire v$RM_11772_out0;
wire v$RM_11773_out0;
wire v$RM_11774_out0;
wire v$RM_11775_out0;
wire v$RM_11776_out0;
wire v$RM_11777_out0;
wire v$RM_11778_out0;
wire v$RM_11779_out0;
wire v$RM_11780_out0;
wire v$RM_11781_out0;
wire v$RM_11782_out0;
wire v$RM_11783_out0;
wire v$RM_11784_out0;
wire v$RM_11785_out0;
wire v$RM_11786_out0;
wire v$RM_11787_out0;
wire v$RM_11788_out0;
wire v$RM_11789_out0;
wire v$RM_11790_out0;
wire v$RM_11791_out0;
wire v$RM_11792_out0;
wire v$RM_11793_out0;
wire v$RM_11794_out0;
wire v$RM_11795_out0;
wire v$RM_11796_out0;
wire v$RM_11797_out0;
wire v$RM_11798_out0;
wire v$RM_11799_out0;
wire v$RM_11800_out0;
wire v$RM_11801_out0;
wire v$RM_11802_out0;
wire v$RM_11803_out0;
wire v$RM_11804_out0;
wire v$RM_11805_out0;
wire v$RM_11806_out0;
wire v$RM_11807_out0;
wire v$RM_11808_out0;
wire v$RM_11809_out0;
wire v$RM_11810_out0;
wire v$RM_11811_out0;
wire v$RM_11812_out0;
wire v$RM_11813_out0;
wire v$RM_11814_out0;
wire v$RM_11815_out0;
wire v$RM_11816_out0;
wire v$RM_11817_out0;
wire v$RM_11818_out0;
wire v$RM_11819_out0;
wire v$RM_11820_out0;
wire v$RM_11821_out0;
wire v$RM_11822_out0;
wire v$RM_11823_out0;
wire v$RM_11824_out0;
wire v$RM_11825_out0;
wire v$RM_11826_out0;
wire v$RM_11827_out0;
wire v$RM_11828_out0;
wire v$RM_11829_out0;
wire v$RM_11830_out0;
wire v$RM_11831_out0;
wire v$RM_11832_out0;
wire v$RM_11833_out0;
wire v$RM_11834_out0;
wire v$RM_11835_out0;
wire v$RM_11836_out0;
wire v$RM_11837_out0;
wire v$RM_11838_out0;
wire v$RM_11839_out0;
wire v$RM_11840_out0;
wire v$RM_11841_out0;
wire v$RM_11842_out0;
wire v$RM_11843_out0;
wire v$RM_11844_out0;
wire v$RM_11845_out0;
wire v$RM_11846_out0;
wire v$RM_11847_out0;
wire v$RM_11848_out0;
wire v$RM_11849_out0;
wire v$RM_11850_out0;
wire v$RM_11851_out0;
wire v$RM_11852_out0;
wire v$RM_11853_out0;
wire v$RM_11854_out0;
wire v$RM_11855_out0;
wire v$RM_11856_out0;
wire v$RM_11857_out0;
wire v$RM_11858_out0;
wire v$RM_11859_out0;
wire v$RM_11860_out0;
wire v$RM_11861_out0;
wire v$RM_11862_out0;
wire v$RM_11863_out0;
wire v$RM_11864_out0;
wire v$RM_11865_out0;
wire v$RM_11866_out0;
wire v$RM_11867_out0;
wire v$RM_11868_out0;
wire v$RM_11869_out0;
wire v$RM_11870_out0;
wire v$RM_11871_out0;
wire v$RM_11872_out0;
wire v$RM_11873_out0;
wire v$RM_11874_out0;
wire v$RM_11875_out0;
wire v$RM_11876_out0;
wire v$RM_11877_out0;
wire v$RM_11878_out0;
wire v$RM_11879_out0;
wire v$RM_11880_out0;
wire v$RM_11881_out0;
wire v$RM_11882_out0;
wire v$RM_11883_out0;
wire v$RM_11884_out0;
wire v$RM_11885_out0;
wire v$RM_11886_out0;
wire v$RM_11887_out0;
wire v$RM_11888_out0;
wire v$RM_11889_out0;
wire v$RM_11890_out0;
wire v$RM_11891_out0;
wire v$RM_11892_out0;
wire v$RM_11893_out0;
wire v$RM_11894_out0;
wire v$RM_11895_out0;
wire v$RM_11896_out0;
wire v$RM_11897_out0;
wire v$RM_11898_out0;
wire v$RM_11899_out0;
wire v$RM_11900_out0;
wire v$RM_11901_out0;
wire v$RM_11902_out0;
wire v$RM_11903_out0;
wire v$RM_11904_out0;
wire v$RM_11905_out0;
wire v$RM_11906_out0;
wire v$RM_11907_out0;
wire v$RM_11908_out0;
wire v$RM_11909_out0;
wire v$RM_11910_out0;
wire v$RM_11911_out0;
wire v$RM_11912_out0;
wire v$RM_11913_out0;
wire v$RM_11914_out0;
wire v$RM_11915_out0;
wire v$RM_11916_out0;
wire v$RM_11917_out0;
wire v$RM_11918_out0;
wire v$RM_11919_out0;
wire v$RM_11920_out0;
wire v$RM_11921_out0;
wire v$RM_11922_out0;
wire v$RM_11923_out0;
wire v$RM_11924_out0;
wire v$RM_11925_out0;
wire v$RM_11926_out0;
wire v$RM_11927_out0;
wire v$RM_11928_out0;
wire v$RM_11929_out0;
wire v$RM_11930_out0;
wire v$RM_11931_out0;
wire v$RM_11932_out0;
wire v$RM_11933_out0;
wire v$RM_11934_out0;
wire v$RM_11935_out0;
wire v$RM_11936_out0;
wire v$RM_11937_out0;
wire v$RM_11938_out0;
wire v$RM_11939_out0;
wire v$RM_11940_out0;
wire v$RM_11941_out0;
wire v$RM_11942_out0;
wire v$RM_11943_out0;
wire v$RM_11944_out0;
wire v$RM_11945_out0;
wire v$RM_11946_out0;
wire v$RM_11947_out0;
wire v$RM_11948_out0;
wire v$RM_11949_out0;
wire v$RM_11950_out0;
wire v$RM_11951_out0;
wire v$RM_11952_out0;
wire v$RM_11953_out0;
wire v$RM_11954_out0;
wire v$RM_11955_out0;
wire v$RM_11956_out0;
wire v$RM_11957_out0;
wire v$RM_11958_out0;
wire v$RM_11959_out0;
wire v$RM_11960_out0;
wire v$RM_11961_out0;
wire v$RM_11962_out0;
wire v$RM_11963_out0;
wire v$RM_11964_out0;
wire v$RM_11965_out0;
wire v$RM_11966_out0;
wire v$RM_11967_out0;
wire v$RM_11968_out0;
wire v$RM_11969_out0;
wire v$RM_11970_out0;
wire v$RM_11971_out0;
wire v$RM_11972_out0;
wire v$RM_11973_out0;
wire v$RM_11974_out0;
wire v$RM_11975_out0;
wire v$RM_11976_out0;
wire v$RM_11977_out0;
wire v$RM_11978_out0;
wire v$RM_11979_out0;
wire v$RM_11980_out0;
wire v$RM_11981_out0;
wire v$RM_11982_out0;
wire v$RM_11983_out0;
wire v$RM_11984_out0;
wire v$RM_11985_out0;
wire v$RM_11986_out0;
wire v$RM_11987_out0;
wire v$RM_11988_out0;
wire v$RM_11989_out0;
wire v$RM_11990_out0;
wire v$RM_11991_out0;
wire v$RM_11992_out0;
wire v$RM_11993_out0;
wire v$RM_11994_out0;
wire v$RM_11995_out0;
wire v$RM_11996_out0;
wire v$RM_11997_out0;
wire v$RM_11998_out0;
wire v$RM_11999_out0;
wire v$RM_12000_out0;
wire v$RM_12001_out0;
wire v$RM_12002_out0;
wire v$RM_12003_out0;
wire v$RM_12004_out0;
wire v$RM_12005_out0;
wire v$RM_12006_out0;
wire v$RM_12007_out0;
wire v$RM_12008_out0;
wire v$RM_12009_out0;
wire v$RM_12010_out0;
wire v$RM_12011_out0;
wire v$RM_12012_out0;
wire v$RM_12013_out0;
wire v$RM_12014_out0;
wire v$RM_12015_out0;
wire v$RM_12016_out0;
wire v$RM_12017_out0;
wire v$RM_12018_out0;
wire v$RM_12019_out0;
wire v$RM_12020_out0;
wire v$RM_12021_out0;
wire v$RM_12022_out0;
wire v$RM_12023_out0;
wire v$RM_12024_out0;
wire v$RM_12025_out0;
wire v$RM_12026_out0;
wire v$RM_12027_out0;
wire v$RM_12028_out0;
wire v$RM_12029_out0;
wire v$RM_12030_out0;
wire v$RM_12031_out0;
wire v$RM_12032_out0;
wire v$RM_12033_out0;
wire v$RM_12034_out0;
wire v$RM_12035_out0;
wire v$RM_12036_out0;
wire v$RM_12037_out0;
wire v$RM_12038_out0;
wire v$RM_12039_out0;
wire v$RM_12040_out0;
wire v$RM_12041_out0;
wire v$RM_12042_out0;
wire v$RM_12043_out0;
wire v$RM_12044_out0;
wire v$RM_12045_out0;
wire v$RM_12046_out0;
wire v$RM_12047_out0;
wire v$RM_12048_out0;
wire v$RM_12049_out0;
wire v$RM_12050_out0;
wire v$RM_12051_out0;
wire v$RM_12052_out0;
wire v$RM_12053_out0;
wire v$RM_12054_out0;
wire v$RM_12055_out0;
wire v$RM_12056_out0;
wire v$RM_12057_out0;
wire v$RM_12058_out0;
wire v$RM_12059_out0;
wire v$RM_12060_out0;
wire v$RM_12061_out0;
wire v$RM_12062_out0;
wire v$RM_12063_out0;
wire v$RM_12064_out0;
wire v$RM_12065_out0;
wire v$RM_12066_out0;
wire v$RM_12067_out0;
wire v$RM_12068_out0;
wire v$RM_12069_out0;
wire v$RM_12070_out0;
wire v$RM_12071_out0;
wire v$RM_12072_out0;
wire v$RM_12073_out0;
wire v$RM_12074_out0;
wire v$RM_12075_out0;
wire v$RM_12076_out0;
wire v$RM_12077_out0;
wire v$RM_12078_out0;
wire v$RM_12079_out0;
wire v$RM_12080_out0;
wire v$RM_12081_out0;
wire v$RM_12082_out0;
wire v$RM_12083_out0;
wire v$RM_12084_out0;
wire v$RM_12085_out0;
wire v$RM_12086_out0;
wire v$RM_12087_out0;
wire v$RM_12088_out0;
wire v$RM_12089_out0;
wire v$RM_12090_out0;
wire v$RM_12091_out0;
wire v$RM_12092_out0;
wire v$RM_12093_out0;
wire v$RM_12094_out0;
wire v$RM_12095_out0;
wire v$RM_12096_out0;
wire v$RM_12097_out0;
wire v$RM_12098_out0;
wire v$RM_12099_out0;
wire v$RM_12100_out0;
wire v$RM_12101_out0;
wire v$RM_12102_out0;
wire v$RM_12103_out0;
wire v$RM_12104_out0;
wire v$RM_12105_out0;
wire v$RM_12106_out0;
wire v$RM_12107_out0;
wire v$RM_12108_out0;
wire v$RM_12109_out0;
wire v$RM_12110_out0;
wire v$RM_12111_out0;
wire v$RM_12112_out0;
wire v$RM_12113_out0;
wire v$RM_12114_out0;
wire v$RM_12115_out0;
wire v$RM_12116_out0;
wire v$RM_12117_out0;
wire v$RM_12118_out0;
wire v$RM_12119_out0;
wire v$RM_12120_out0;
wire v$RM_12121_out0;
wire v$RM_12122_out0;
wire v$RM_12123_out0;
wire v$RM_12124_out0;
wire v$RM_12125_out0;
wire v$RM_12126_out0;
wire v$RM_12127_out0;
wire v$RM_12128_out0;
wire v$RM_12129_out0;
wire v$RM_12130_out0;
wire v$RM_12131_out0;
wire v$RM_12132_out0;
wire v$RM_12133_out0;
wire v$RM_12134_out0;
wire v$RM_12135_out0;
wire v$RM_12136_out0;
wire v$RM_12137_out0;
wire v$RM_12138_out0;
wire v$RM_12139_out0;
wire v$RM_12140_out0;
wire v$RM_12141_out0;
wire v$RM_12142_out0;
wire v$RM_12143_out0;
wire v$RM_12144_out0;
wire v$RM_12145_out0;
wire v$RM_12146_out0;
wire v$RM_12147_out0;
wire v$RM_12148_out0;
wire v$RM_12149_out0;
wire v$RM_12150_out0;
wire v$RM_12151_out0;
wire v$RM_12152_out0;
wire v$RM_12153_out0;
wire v$RM_12154_out0;
wire v$RM_12155_out0;
wire v$RM_12156_out0;
wire v$RM_12157_out0;
wire v$RM_12158_out0;
wire v$RM_12159_out0;
wire v$RM_12160_out0;
wire v$RM_12161_out0;
wire v$RM_12162_out0;
wire v$RM_12163_out0;
wire v$RM_12164_out0;
wire v$RM_12165_out0;
wire v$RM_12166_out0;
wire v$RM_12167_out0;
wire v$RM_12168_out0;
wire v$RM_12169_out0;
wire v$RM_12170_out0;
wire v$RM_12171_out0;
wire v$RM_12172_out0;
wire v$RM_12173_out0;
wire v$RM_12174_out0;
wire v$RM_12175_out0;
wire v$RM_12176_out0;
wire v$RM_12177_out0;
wire v$RM_12178_out0;
wire v$RM_12179_out0;
wire v$RM_12180_out0;
wire v$RM_12181_out0;
wire v$RM_12182_out0;
wire v$RM_12183_out0;
wire v$RM_12184_out0;
wire v$RM_12185_out0;
wire v$RM_12186_out0;
wire v$RM_12187_out0;
wire v$RM_12188_out0;
wire v$RM_12189_out0;
wire v$RM_12190_out0;
wire v$RM_12191_out0;
wire v$RM_12192_out0;
wire v$RM_12193_out0;
wire v$RM_12194_out0;
wire v$RM_12195_out0;
wire v$RM_12196_out0;
wire v$RM_12197_out0;
wire v$RM_12198_out0;
wire v$RM_12199_out0;
wire v$RM_12200_out0;
wire v$RM_12201_out0;
wire v$RM_12202_out0;
wire v$RM_12203_out0;
wire v$RM_12204_out0;
wire v$RM_12205_out0;
wire v$RM_12206_out0;
wire v$RM_12207_out0;
wire v$RM_12208_out0;
wire v$RM_12209_out0;
wire v$RM_12210_out0;
wire v$RM_12211_out0;
wire v$RM_12212_out0;
wire v$RM_12213_out0;
wire v$RM_12214_out0;
wire v$RM_12215_out0;
wire v$RM_12216_out0;
wire v$RM_12217_out0;
wire v$RM_12218_out0;
wire v$RM_12219_out0;
wire v$RM_12220_out0;
wire v$RM_12221_out0;
wire v$RM_12222_out0;
wire v$RM_12223_out0;
wire v$RM_12224_out0;
wire v$RM_12225_out0;
wire v$RM_12226_out0;
wire v$RM_12227_out0;
wire v$RM_12228_out0;
wire v$RM_12229_out0;
wire v$RM_3355_out0;
wire v$RM_3356_out0;
wire v$RM_3357_out0;
wire v$RM_3358_out0;
wire v$RM_3359_out0;
wire v$RM_3360_out0;
wire v$RM_3361_out0;
wire v$RM_3362_out0;
wire v$RM_3363_out0;
wire v$RM_3364_out0;
wire v$RM_3365_out0;
wire v$RM_3366_out0;
wire v$RM_3367_out0;
wire v$RM_3368_out0;
wire v$RM_3369_out0;
wire v$RM_3370_out0;
wire v$RM_3371_out0;
wire v$RM_3372_out0;
wire v$RM_3373_out0;
wire v$RM_3374_out0;
wire v$RM_3375_out0;
wire v$RM_3376_out0;
wire v$RM_3377_out0;
wire v$RM_3378_out0;
wire v$RM_3379_out0;
wire v$RM_3380_out0;
wire v$RM_3381_out0;
wire v$RM_3382_out0;
wire v$RM_3383_out0;
wire v$RM_3384_out0;
wire v$RM_3385_out0;
wire v$RM_3386_out0;
wire v$RM_3387_out0;
wire v$RM_3388_out0;
wire v$RM_3389_out0;
wire v$RM_3390_out0;
wire v$RM_3391_out0;
wire v$RM_3392_out0;
wire v$RM_3393_out0;
wire v$RM_3394_out0;
wire v$RM_3395_out0;
wire v$RM_3396_out0;
wire v$RM_3397_out0;
wire v$RM_3398_out0;
wire v$RM_3399_out0;
wire v$RM_3400_out0;
wire v$RM_3401_out0;
wire v$RM_3402_out0;
wire v$RM_3403_out0;
wire v$RM_3404_out0;
wire v$RM_3405_out0;
wire v$RM_3406_out0;
wire v$RM_3407_out0;
wire v$RM_3408_out0;
wire v$RM_3409_out0;
wire v$RM_3410_out0;
wire v$RM_3411_out0;
wire v$RM_3412_out0;
wire v$RM_3413_out0;
wire v$RM_3414_out0;
wire v$RM_3415_out0;
wire v$RM_3416_out0;
wire v$RM_3417_out0;
wire v$RM_3418_out0;
wire v$RM_3419_out0;
wire v$RM_3420_out0;
wire v$RM_3421_out0;
wire v$RM_3422_out0;
wire v$RM_3423_out0;
wire v$RM_3424_out0;
wire v$RM_3425_out0;
wire v$RM_3426_out0;
wire v$RM_3427_out0;
wire v$RM_3428_out0;
wire v$RM_3429_out0;
wire v$RM_3430_out0;
wire v$RM_3431_out0;
wire v$RM_3432_out0;
wire v$RM_3433_out0;
wire v$RM_3434_out0;
wire v$RM_3435_out0;
wire v$RM_3436_out0;
wire v$RM_3437_out0;
wire v$RM_3438_out0;
wire v$RM_3439_out0;
wire v$RM_3440_out0;
wire v$RM_3441_out0;
wire v$RM_3442_out0;
wire v$RM_3443_out0;
wire v$RM_3444_out0;
wire v$RM_3445_out0;
wire v$RM_3446_out0;
wire v$RM_3447_out0;
wire v$RM_3448_out0;
wire v$RM_3449_out0;
wire v$RM_3450_out0;
wire v$RM_3451_out0;
wire v$RM_3452_out0;
wire v$RM_3453_out0;
wire v$RM_3454_out0;
wire v$RM_3455_out0;
wire v$RM_3456_out0;
wire v$RM_3457_out0;
wire v$RM_3458_out0;
wire v$RM_3459_out0;
wire v$RM_3460_out0;
wire v$RM_3461_out0;
wire v$RM_3462_out0;
wire v$RM_3463_out0;
wire v$RM_3464_out0;
wire v$RM_3465_out0;
wire v$RM_3466_out0;
wire v$RM_3467_out0;
wire v$RM_3468_out0;
wire v$RM_3469_out0;
wire v$RM_3470_out0;
wire v$RM_3471_out0;
wire v$RM_3472_out0;
wire v$RM_3473_out0;
wire v$RM_3474_out0;
wire v$RM_3475_out0;
wire v$RM_3476_out0;
wire v$RM_3477_out0;
wire v$RM_3478_out0;
wire v$RM_3479_out0;
wire v$RM_3480_out0;
wire v$RM_3481_out0;
wire v$RM_3482_out0;
wire v$RM_3483_out0;
wire v$RM_3484_out0;
wire v$RM_3485_out0;
wire v$RM_3486_out0;
wire v$RM_3487_out0;
wire v$RM_3488_out0;
wire v$RM_3489_out0;
wire v$RM_3490_out0;
wire v$RM_3491_out0;
wire v$RM_3492_out0;
wire v$RM_3493_out0;
wire v$RM_3494_out0;
wire v$RM_3495_out0;
wire v$RM_3496_out0;
wire v$RM_3497_out0;
wire v$RM_3498_out0;
wire v$RM_3499_out0;
wire v$RM_3500_out0;
wire v$RM_3501_out0;
wire v$RM_3502_out0;
wire v$RM_3503_out0;
wire v$RM_3504_out0;
wire v$RM_3505_out0;
wire v$RM_3506_out0;
wire v$RM_3507_out0;
wire v$RM_3508_out0;
wire v$RM_3509_out0;
wire v$RM_3510_out0;
wire v$RM_3511_out0;
wire v$RM_3512_out0;
wire v$RM_3513_out0;
wire v$RM_3514_out0;
wire v$RM_3515_out0;
wire v$RM_3516_out0;
wire v$RM_3517_out0;
wire v$RM_3518_out0;
wire v$RM_3519_out0;
wire v$RM_3520_out0;
wire v$RM_3521_out0;
wire v$RM_3522_out0;
wire v$RM_3523_out0;
wire v$RM_3524_out0;
wire v$RM_3525_out0;
wire v$RM_3526_out0;
wire v$RM_3527_out0;
wire v$RM_3528_out0;
wire v$RM_3529_out0;
wire v$RM_3530_out0;
wire v$RM_3531_out0;
wire v$RM_3532_out0;
wire v$RM_3533_out0;
wire v$RM_3534_out0;
wire v$RM_3535_out0;
wire v$RM_3536_out0;
wire v$RM_3537_out0;
wire v$RM_3538_out0;
wire v$RM_3539_out0;
wire v$RM_3540_out0;
wire v$RM_3541_out0;
wire v$RM_3542_out0;
wire v$RM_3543_out0;
wire v$RM_3544_out0;
wire v$RM_3545_out0;
wire v$RM_3546_out0;
wire v$RM_3547_out0;
wire v$RM_3548_out0;
wire v$RM_3549_out0;
wire v$RM_3550_out0;
wire v$RM_3551_out0;
wire v$RM_3552_out0;
wire v$RM_3553_out0;
wire v$RM_3554_out0;
wire v$RM_3555_out0;
wire v$RM_3556_out0;
wire v$RM_3557_out0;
wire v$RM_3558_out0;
wire v$RM_3559_out0;
wire v$RM_3560_out0;
wire v$RM_3561_out0;
wire v$RM_3562_out0;
wire v$RM_3563_out0;
wire v$RM_3564_out0;
wire v$RM_3565_out0;
wire v$RM_3566_out0;
wire v$RM_3567_out0;
wire v$RM_3568_out0;
wire v$RM_3569_out0;
wire v$RM_3570_out0;
wire v$RM_3571_out0;
wire v$RM_3572_out0;
wire v$RM_3573_out0;
wire v$RM_3574_out0;
wire v$RM_3575_out0;
wire v$RM_3576_out0;
wire v$RM_3577_out0;
wire v$RM_3578_out0;
wire v$RM_3579_out0;
wire v$RM_3580_out0;
wire v$RM_3581_out0;
wire v$RM_3582_out0;
wire v$RM_3583_out0;
wire v$RM_3584_out0;
wire v$RM_3585_out0;
wire v$RM_3586_out0;
wire v$RM_3587_out0;
wire v$RM_3588_out0;
wire v$RM_3589_out0;
wire v$RM_3590_out0;
wire v$RM_3591_out0;
wire v$RM_3592_out0;
wire v$RM_3593_out0;
wire v$RM_3594_out0;
wire v$RM_3595_out0;
wire v$RM_3596_out0;
wire v$RM_3597_out0;
wire v$RM_3598_out0;
wire v$RM_3599_out0;
wire v$RM_3600_out0;
wire v$RM_3601_out0;
wire v$RM_3602_out0;
wire v$RM_3603_out0;
wire v$RM_3604_out0;
wire v$RM_3605_out0;
wire v$RM_3606_out0;
wire v$RM_3607_out0;
wire v$RM_3608_out0;
wire v$RM_3609_out0;
wire v$RM_3610_out0;
wire v$RM_3611_out0;
wire v$RM_3612_out0;
wire v$RM_3613_out0;
wire v$RM_3614_out0;
wire v$RM_3615_out0;
wire v$RM_3616_out0;
wire v$RM_3617_out0;
wire v$RM_3618_out0;
wire v$RM_3619_out0;
wire v$RM_3620_out0;
wire v$RM_3621_out0;
wire v$RM_3622_out0;
wire v$RM_3623_out0;
wire v$RM_3624_out0;
wire v$RM_3625_out0;
wire v$RM_3626_out0;
wire v$RM_3627_out0;
wire v$RM_3628_out0;
wire v$RM_3629_out0;
wire v$RM_3630_out0;
wire v$RM_3631_out0;
wire v$RM_3632_out0;
wire v$RM_3633_out0;
wire v$RM_3634_out0;
wire v$RM_3635_out0;
wire v$RM_3636_out0;
wire v$RM_3637_out0;
wire v$RM_3638_out0;
wire v$RM_3639_out0;
wire v$RM_3640_out0;
wire v$RM_3641_out0;
wire v$RM_3642_out0;
wire v$RM_3643_out0;
wire v$RM_3644_out0;
wire v$RM_3645_out0;
wire v$RM_3646_out0;
wire v$RM_3647_out0;
wire v$RM_3648_out0;
wire v$RM_3649_out0;
wire v$RM_3650_out0;
wire v$RM_3651_out0;
wire v$RM_3652_out0;
wire v$RM_3653_out0;
wire v$RM_3654_out0;
wire v$RM_3655_out0;
wire v$RM_3656_out0;
wire v$RM_3657_out0;
wire v$RM_3658_out0;
wire v$RM_3659_out0;
wire v$RM_3660_out0;
wire v$RM_3661_out0;
wire v$RM_3662_out0;
wire v$RM_3663_out0;
wire v$RM_3664_out0;
wire v$RM_3665_out0;
wire v$RM_3666_out0;
wire v$RM_3667_out0;
wire v$RM_3668_out0;
wire v$RM_3669_out0;
wire v$RM_3670_out0;
wire v$RM_3671_out0;
wire v$RM_3672_out0;
wire v$RM_3673_out0;
wire v$RM_3674_out0;
wire v$RM_3675_out0;
wire v$RM_3676_out0;
wire v$RM_3677_out0;
wire v$RM_3678_out0;
wire v$RM_3679_out0;
wire v$RM_3680_out0;
wire v$RM_3681_out0;
wire v$RM_3682_out0;
wire v$RM_3683_out0;
wire v$RM_3684_out0;
wire v$RM_3685_out0;
wire v$RM_3686_out0;
wire v$RM_3687_out0;
wire v$RM_3688_out0;
wire v$RM_3689_out0;
wire v$RM_3690_out0;
wire v$RM_3691_out0;
wire v$RM_3692_out0;
wire v$RM_3693_out0;
wire v$RM_3694_out0;
wire v$RM_3695_out0;
wire v$RM_3696_out0;
wire v$RM_3697_out0;
wire v$RM_3698_out0;
wire v$RM_3699_out0;
wire v$RM_3700_out0;
wire v$RM_3701_out0;
wire v$RM_3702_out0;
wire v$RM_3703_out0;
wire v$RM_3704_out0;
wire v$RM_3705_out0;
wire v$RM_3706_out0;
wire v$RM_3707_out0;
wire v$RM_3708_out0;
wire v$RM_3709_out0;
wire v$RM_3710_out0;
wire v$RM_3711_out0;
wire v$RM_3712_out0;
wire v$RM_3713_out0;
wire v$RM_3714_out0;
wire v$RM_3715_out0;
wire v$RM_3716_out0;
wire v$RM_3717_out0;
wire v$RM_3718_out0;
wire v$RM_3719_out0;
wire v$RM_3720_out0;
wire v$RM_3721_out0;
wire v$RM_3722_out0;
wire v$RM_3723_out0;
wire v$RM_3724_out0;
wire v$RM_3725_out0;
wire v$RM_3726_out0;
wire v$RM_3727_out0;
wire v$RM_3728_out0;
wire v$RM_3729_out0;
wire v$RM_3730_out0;
wire v$RM_3731_out0;
wire v$RM_3732_out0;
wire v$RM_3733_out0;
wire v$RM_3734_out0;
wire v$RM_3735_out0;
wire v$RM_3736_out0;
wire v$RM_3737_out0;
wire v$RM_3738_out0;
wire v$RM_3739_out0;
wire v$RM_3740_out0;
wire v$RM_3741_out0;
wire v$RM_3742_out0;
wire v$RM_3743_out0;
wire v$RM_3744_out0;
wire v$RM_3745_out0;
wire v$RM_3746_out0;
wire v$RM_3747_out0;
wire v$RM_3748_out0;
wire v$RM_3749_out0;
wire v$RM_3750_out0;
wire v$RM_3751_out0;
wire v$RM_3752_out0;
wire v$RM_3753_out0;
wire v$RM_3754_out0;
wire v$RM_3755_out0;
wire v$RM_3756_out0;
wire v$RM_3757_out0;
wire v$RM_3758_out0;
wire v$RM_3759_out0;
wire v$RM_3760_out0;
wire v$RM_3761_out0;
wire v$RM_3762_out0;
wire v$RM_3763_out0;
wire v$RM_3764_out0;
wire v$RM_3765_out0;
wire v$RM_3766_out0;
wire v$RM_3767_out0;
wire v$RM_3768_out0;
wire v$RM_3769_out0;
wire v$RM_3770_out0;
wire v$RM_3771_out0;
wire v$RM_3772_out0;
wire v$RM_3773_out0;
wire v$RM_3774_out0;
wire v$RM_3775_out0;
wire v$RM_3776_out0;
wire v$RM_3777_out0;
wire v$RM_3778_out0;
wire v$RM_3779_out0;
wire v$RM_3780_out0;
wire v$RM_3781_out0;
wire v$RM_3782_out0;
wire v$RM_3783_out0;
wire v$RM_3784_out0;
wire v$RM_3785_out0;
wire v$RM_3786_out0;
wire v$RM_3787_out0;
wire v$RM_3788_out0;
wire v$RM_3789_out0;
wire v$RM_3790_out0;
wire v$RM_3791_out0;
wire v$RM_3792_out0;
wire v$RM_3793_out0;
wire v$RM_3794_out0;
wire v$RM_3795_out0;
wire v$RM_3796_out0;
wire v$RM_3797_out0;
wire v$RM_3798_out0;
wire v$RM_3799_out0;
wire v$RM_3800_out0;
wire v$RM_3801_out0;
wire v$RM_3802_out0;
wire v$ROM1_462_out0;
wire v$ROR_282_out0;
wire v$ROR_283_out0;
wire v$ROR_3286_out0;
wire v$ROR_3287_out0;
wire v$ROR_3288_out0;
wire v$ROR_3289_out0;
wire v$ROR_544_out0;
wire v$ROR_545_out0;
wire v$RX$BYTE$READY_2436_out0;
wire v$RX$BYTEREADY_8756_out0;
wire v$RX$DONE$RECEIVING_10484_out0;
wire v$RX$INST0_2970_out0;
wire v$RX$INST1_12_out0;
wire v$RX$INSTRUCTION_11170_out0;
wire v$RX$INSTRUCTION_11171_out0;
wire v$RX$INSTRUCTION_13325_out0;
wire v$RX$INSTRUCTION_2343_out0;
wire v$RX$INSTRUCTION_2344_out0;
wire v$RX$INSTRUCTION_3258_out0;
wire v$RX$INSTRUCTION_3259_out0;
wire v$RX$INSTRUCTION_4659_out0;
wire v$RX$INSTRUCTION_8686_out0;
wire v$RX$INSTRUCTION_94_out0;
wire v$RX$INSTRUCTION_95_out0;
wire v$RX$INST_2334_out0;
wire v$RX$OVERFLOW_426_out0;
wire v$RX$OVERFLOW_4469_out0;
wire v$RX$OVERFLOW_5848_out0;
wire v$RXBYTERECEIVED_3269_out0;
wire v$RXBYTERECEIVED_91_out0;
wire v$SBC_11051_out0;
wire v$SBC_11052_out0;
wire v$SBC_13605_out0;
wire v$SBC_13606_out0;
wire v$SBC_4825_out0;
wire v$SBC_4826_out0;
wire v$SEL1_10304_out0;
wire v$SEL1_1164_out0;
wire v$SEL1_1204_out0;
wire v$SEL1_13445_out0;
wire v$SEL1_2305_out0;
wire v$SEL1_2306_out0;
wire v$SEL1_2319_out0;
wire v$SEL1_240_out0;
wire v$SEL1_2428_out0;
wire v$SEL1_2914_out0;
wire v$SEL1_2915_out0;
wire v$SEL1_4858_out0;
wire v$SEL2_10323_out0;
wire v$SEL2_10324_out0;
wire v$SEL2_280_out0;
wire v$SEL2_281_out0;
wire v$SEL3_1143_out0;
wire v$SEL3_1144_out0;
wire v$SEL3_2615_out0;
wire v$SEL3_2616_out0;
wire v$SEL4_7636_out0;
wire v$SEL4_7637_out0;
wire v$SEL5_3049_out0;
wire v$SEL5_3050_out0;
wire v$SHIFHT$ENABLE_13500_out0;
wire v$SHIFHT$ENABLE_13501_out0;
wire v$SHIFHT$ENABLE_13502_out0;
wire v$SHIFHT$ENABLE_13503_out0;
wire v$SHIFT$ENABLE_8684_out0;
wire v$SHIFT$RD_2544_out0;
wire v$SHIFT$RD_2545_out0;
wire v$SHIFT$WHICH$OP_10465_out0;
wire v$SHIFT$WHICH$OP_10466_out0;
wire v$SHIFT$WHICH$OP_10715_out0;
wire v$SHIFT$WHICH$OP_10716_out0;
wire v$SHIFT$WHICH$OP_4459_out0;
wire v$SHIFT$WHICH$OP_4460_out0;
wire v$SIGN$ANS_10302_out0;
wire v$SIGN$ANS_10303_out0;
wire v$SIGN$ANS_1970_out0;
wire v$SIGN$ANS_1971_out0;
wire v$SIGN$ANS_4457_out0;
wire v$SIGN$ANS_4458_out0;
wire v$SIGN$ANS_8650_out0;
wire v$SIGN$ANS_8651_out0;
wire v$STALL$DUAL$CORE_12234_out0;
wire v$STALL$DUAL$CORE_12235_out0;
wire v$STALL$DUAL$CORE_13617_out0;
wire v$STALL$DUAL$CORE_13618_out0;
wire v$STALL$DUAL$CORE_1738_out0;
wire v$STALL$DUAL$CORE_1739_out0;
wire v$STALL$DUAL$CORE_1958_out0;
wire v$STALL$DUAL$CORE_1959_out0;
wire v$STALL$DUAL$CORE_3127_out0;
wire v$STALL$DUAL$CORE_3128_out0;
wire v$STALL$DUAL$CORE_3264_out0;
wire v$STALL$DUAL$CORE_3265_out0;
wire v$STALL$DUAL$CORE_4695_out0;
wire v$STALL$DUAL$CORE_4696_out0;
wire v$STALL$dual$core_8741_out0;
wire v$STALL$dual$core_8742_out0;
wire v$STALL_10281_out0;
wire v$STALL_10282_out0;
wire v$STALL_1758_out0;
wire v$STALL_1759_out0;
wire v$STALL_427_out0;
wire v$STALL_428_out0;
wire v$STALL_6910_out0;
wire v$STALL_6911_out0;
wire v$STARTBIT_6967_out0;
wire v$STARTBIT_6968_out0;
wire v$STARTBIT_6969_out0;
wire v$STARTBIT_6970_out0;
wire v$START_13394_out0;
wire v$START_13395_out0;
wire v$START_3027_out0;
wire v$START_3028_out0;
wire v$START_392_out0;
wire v$START_393_out0;
wire v$STAT$INSTRUCTION_10272_out0;
wire v$STAT$INSTRUCTION_10273_out0;
wire v$STAT$INSTRUCTION_2434_out0;
wire v$STAT$INSTRUCTION_2435_out0;
wire v$STAT$INSTRUCTION_2855_out0;
wire v$STAT$INSTRUCTION_2856_out0;
wire v$STORE$PCOUNTER_2102_out0;
wire v$STORE$PCOUNTER_2103_out0;
wire v$STORE$WEN_4544_out0;
wire v$STORE$WEN_4545_out0;
wire v$STORE$pccounter_2883_out0;
wire v$STORE$pccounter_2884_out0;
wire v$STORE_10831_out0;
wire v$STORE_10832_out0;
wire v$STORE_1195_out0;
wire v$STORE_1196_out0;
wire v$STORE_12245_out0;
wire v$STORE_12246_out0;
wire v$STORE_13298_out0;
wire v$STORE_13299_out0;
wire v$STORE_221_out0;
wire v$STORE_222_out0;
wire v$STORE_540_out0;
wire v$STORE_541_out0;
wire v$STP_10307_out0;
wire v$STP_10308_out0;
wire v$STP_10352_out0;
wire v$STP_10353_out0;
wire v$STP_10467_out0;
wire v$STP_10468_out0;
wire v$STP_10977_out0;
wire v$STP_10978_out0;
wire v$STP_11240_out0;
wire v$STP_11241_out0;
wire v$STP_52_out0;
wire v$STP_53_out0;
wire v$SUB$INSTRUCTION_11195_out0;
wire v$SUB$INSTRUCTION_11196_out0;
wire v$SUB$INSTRUCTION_2789_out0;
wire v$SUB$INSTRUCTION_2790_out0;
wire v$SUB$INSTRUCTION_7085_out0;
wire v$SUB$INSTRUCTION_7086_out0;
wire v$SUBNORMAL_8808_out0;
wire v$SUBNORMAL_8809_out0;
wire v$SUB_12247_out0;
wire v$SUB_12248_out0;
wire v$SUB_2695_out0;
wire v$SUB_2696_out0;
wire v$SUB_2909_out0;
wire v$SUB_2910_out0;
wire v$SUB_2957_out0;
wire v$SUB_2958_out0;
wire v$SUB_4616_out0;
wire v$SUB_4617_out0;
wire v$SUB_4618_out0;
wire v$SUB_4619_out0;
wire v$SUB_8663_out0;
wire v$SUB_8664_out0;
wire v$S_11300_out0;
wire v$S_11301_out0;
wire v$S_1219_out0;
wire v$S_1220_out0;
wire v$S_1221_out0;
wire v$S_1222_out0;
wire v$S_1223_out0;
wire v$S_1224_out0;
wire v$S_1225_out0;
wire v$S_1226_out0;
wire v$S_1227_out0;
wire v$S_1228_out0;
wire v$S_1229_out0;
wire v$S_1230_out0;
wire v$S_1231_out0;
wire v$S_1232_out0;
wire v$S_1233_out0;
wire v$S_1234_out0;
wire v$S_1235_out0;
wire v$S_1236_out0;
wire v$S_1237_out0;
wire v$S_1238_out0;
wire v$S_1239_out0;
wire v$S_1240_out0;
wire v$S_1241_out0;
wire v$S_1242_out0;
wire v$S_1243_out0;
wire v$S_1244_out0;
wire v$S_1245_out0;
wire v$S_1246_out0;
wire v$S_1247_out0;
wire v$S_1248_out0;
wire v$S_1249_out0;
wire v$S_1250_out0;
wire v$S_1251_out0;
wire v$S_1252_out0;
wire v$S_1253_out0;
wire v$S_1254_out0;
wire v$S_1255_out0;
wire v$S_1256_out0;
wire v$S_1257_out0;
wire v$S_1258_out0;
wire v$S_1259_out0;
wire v$S_1260_out0;
wire v$S_1261_out0;
wire v$S_1262_out0;
wire v$S_1263_out0;
wire v$S_1264_out0;
wire v$S_1265_out0;
wire v$S_1266_out0;
wire v$S_1267_out0;
wire v$S_1268_out0;
wire v$S_1269_out0;
wire v$S_1270_out0;
wire v$S_1271_out0;
wire v$S_1272_out0;
wire v$S_1273_out0;
wire v$S_1274_out0;
wire v$S_1275_out0;
wire v$S_1276_out0;
wire v$S_1277_out0;
wire v$S_1278_out0;
wire v$S_1279_out0;
wire v$S_1280_out0;
wire v$S_1281_out0;
wire v$S_1282_out0;
wire v$S_1283_out0;
wire v$S_1284_out0;
wire v$S_1285_out0;
wire v$S_1286_out0;
wire v$S_1287_out0;
wire v$S_1288_out0;
wire v$S_1289_out0;
wire v$S_1290_out0;
wire v$S_1291_out0;
wire v$S_1292_out0;
wire v$S_1293_out0;
wire v$S_1294_out0;
wire v$S_1295_out0;
wire v$S_1296_out0;
wire v$S_1297_out0;
wire v$S_1298_out0;
wire v$S_1299_out0;
wire v$S_1300_out0;
wire v$S_1301_out0;
wire v$S_1302_out0;
wire v$S_1303_out0;
wire v$S_1304_out0;
wire v$S_1305_out0;
wire v$S_1306_out0;
wire v$S_1307_out0;
wire v$S_1308_out0;
wire v$S_1309_out0;
wire v$S_1310_out0;
wire v$S_1311_out0;
wire v$S_1312_out0;
wire v$S_1313_out0;
wire v$S_1314_out0;
wire v$S_1315_out0;
wire v$S_1316_out0;
wire v$S_1317_out0;
wire v$S_1318_out0;
wire v$S_1319_out0;
wire v$S_1320_out0;
wire v$S_1321_out0;
wire v$S_1322_out0;
wire v$S_1323_out0;
wire v$S_1324_out0;
wire v$S_1325_out0;
wire v$S_1326_out0;
wire v$S_1327_out0;
wire v$S_1328_out0;
wire v$S_1329_out0;
wire v$S_1330_out0;
wire v$S_1331_out0;
wire v$S_1332_out0;
wire v$S_1333_out0;
wire v$S_1334_out0;
wire v$S_1335_out0;
wire v$S_1336_out0;
wire v$S_1337_out0;
wire v$S_1338_out0;
wire v$S_1339_out0;
wire v$S_1340_out0;
wire v$S_1341_out0;
wire v$S_1342_out0;
wire v$S_1343_out0;
wire v$S_1344_out0;
wire v$S_1345_out0;
wire v$S_1346_out0;
wire v$S_1347_out0;
wire v$S_1348_out0;
wire v$S_1349_out0;
wire v$S_1350_out0;
wire v$S_1351_out0;
wire v$S_1352_out0;
wire v$S_1353_out0;
wire v$S_1354_out0;
wire v$S_1355_out0;
wire v$S_1356_out0;
wire v$S_1357_out0;
wire v$S_1358_out0;
wire v$S_1359_out0;
wire v$S_1360_out0;
wire v$S_1361_out0;
wire v$S_1362_out0;
wire v$S_1363_out0;
wire v$S_1364_out0;
wire v$S_1365_out0;
wire v$S_1366_out0;
wire v$S_1367_out0;
wire v$S_1368_out0;
wire v$S_1369_out0;
wire v$S_1370_out0;
wire v$S_1371_out0;
wire v$S_1372_out0;
wire v$S_1373_out0;
wire v$S_1374_out0;
wire v$S_1375_out0;
wire v$S_1376_out0;
wire v$S_1377_out0;
wire v$S_1378_out0;
wire v$S_1379_out0;
wire v$S_1380_out0;
wire v$S_1381_out0;
wire v$S_1382_out0;
wire v$S_1383_out0;
wire v$S_1384_out0;
wire v$S_1385_out0;
wire v$S_1386_out0;
wire v$S_1387_out0;
wire v$S_1388_out0;
wire v$S_1389_out0;
wire v$S_1390_out0;
wire v$S_1391_out0;
wire v$S_1392_out0;
wire v$S_1393_out0;
wire v$S_1394_out0;
wire v$S_1395_out0;
wire v$S_1396_out0;
wire v$S_1397_out0;
wire v$S_1398_out0;
wire v$S_1399_out0;
wire v$S_1400_out0;
wire v$S_1401_out0;
wire v$S_1402_out0;
wire v$S_1403_out0;
wire v$S_1404_out0;
wire v$S_1405_out0;
wire v$S_1406_out0;
wire v$S_1407_out0;
wire v$S_1408_out0;
wire v$S_1409_out0;
wire v$S_1410_out0;
wire v$S_1411_out0;
wire v$S_1412_out0;
wire v$S_1413_out0;
wire v$S_1414_out0;
wire v$S_1415_out0;
wire v$S_1416_out0;
wire v$S_1417_out0;
wire v$S_1418_out0;
wire v$S_1419_out0;
wire v$S_1420_out0;
wire v$S_1421_out0;
wire v$S_1422_out0;
wire v$S_1423_out0;
wire v$S_1424_out0;
wire v$S_1425_out0;
wire v$S_1426_out0;
wire v$S_1427_out0;
wire v$S_1428_out0;
wire v$S_1429_out0;
wire v$S_1430_out0;
wire v$S_1431_out0;
wire v$S_1432_out0;
wire v$S_1433_out0;
wire v$S_1434_out0;
wire v$S_1435_out0;
wire v$S_1436_out0;
wire v$S_1437_out0;
wire v$S_1438_out0;
wire v$S_1439_out0;
wire v$S_1440_out0;
wire v$S_1441_out0;
wire v$S_1442_out0;
wire v$S_1443_out0;
wire v$S_1444_out0;
wire v$S_1445_out0;
wire v$S_1446_out0;
wire v$S_1447_out0;
wire v$S_1448_out0;
wire v$S_1449_out0;
wire v$S_1450_out0;
wire v$S_1451_out0;
wire v$S_1452_out0;
wire v$S_1453_out0;
wire v$S_1454_out0;
wire v$S_1455_out0;
wire v$S_1456_out0;
wire v$S_1457_out0;
wire v$S_1458_out0;
wire v$S_1459_out0;
wire v$S_1460_out0;
wire v$S_1461_out0;
wire v$S_1462_out0;
wire v$S_1463_out0;
wire v$S_1464_out0;
wire v$S_1465_out0;
wire v$S_1466_out0;
wire v$S_1467_out0;
wire v$S_1468_out0;
wire v$S_1469_out0;
wire v$S_1470_out0;
wire v$S_1471_out0;
wire v$S_1472_out0;
wire v$S_1473_out0;
wire v$S_1474_out0;
wire v$S_1475_out0;
wire v$S_1476_out0;
wire v$S_1477_out0;
wire v$S_1478_out0;
wire v$S_1479_out0;
wire v$S_1480_out0;
wire v$S_1481_out0;
wire v$S_1482_out0;
wire v$S_1483_out0;
wire v$S_1484_out0;
wire v$S_1485_out0;
wire v$S_1486_out0;
wire v$S_1487_out0;
wire v$S_1488_out0;
wire v$S_1489_out0;
wire v$S_1490_out0;
wire v$S_1491_out0;
wire v$S_1492_out0;
wire v$S_1493_out0;
wire v$S_1494_out0;
wire v$S_1495_out0;
wire v$S_1496_out0;
wire v$S_1497_out0;
wire v$S_1498_out0;
wire v$S_1499_out0;
wire v$S_1500_out0;
wire v$S_1501_out0;
wire v$S_1502_out0;
wire v$S_1503_out0;
wire v$S_1504_out0;
wire v$S_1505_out0;
wire v$S_1506_out0;
wire v$S_1507_out0;
wire v$S_1508_out0;
wire v$S_1509_out0;
wire v$S_1510_out0;
wire v$S_1511_out0;
wire v$S_1512_out0;
wire v$S_1513_out0;
wire v$S_1514_out0;
wire v$S_1515_out0;
wire v$S_1516_out0;
wire v$S_1517_out0;
wire v$S_1518_out0;
wire v$S_1519_out0;
wire v$S_1520_out0;
wire v$S_1521_out0;
wire v$S_1522_out0;
wire v$S_1523_out0;
wire v$S_1524_out0;
wire v$S_1525_out0;
wire v$S_1526_out0;
wire v$S_1527_out0;
wire v$S_1528_out0;
wire v$S_1529_out0;
wire v$S_1530_out0;
wire v$S_1531_out0;
wire v$S_1532_out0;
wire v$S_1533_out0;
wire v$S_1534_out0;
wire v$S_1535_out0;
wire v$S_1536_out0;
wire v$S_1537_out0;
wire v$S_1538_out0;
wire v$S_1539_out0;
wire v$S_1540_out0;
wire v$S_1541_out0;
wire v$S_1542_out0;
wire v$S_1543_out0;
wire v$S_1544_out0;
wire v$S_1545_out0;
wire v$S_1546_out0;
wire v$S_1547_out0;
wire v$S_1548_out0;
wire v$S_1549_out0;
wire v$S_1550_out0;
wire v$S_1551_out0;
wire v$S_1552_out0;
wire v$S_1553_out0;
wire v$S_1554_out0;
wire v$S_1555_out0;
wire v$S_1556_out0;
wire v$S_1557_out0;
wire v$S_1558_out0;
wire v$S_1559_out0;
wire v$S_1560_out0;
wire v$S_1561_out0;
wire v$S_1562_out0;
wire v$S_1563_out0;
wire v$S_1564_out0;
wire v$S_1565_out0;
wire v$S_1566_out0;
wire v$S_1567_out0;
wire v$S_1568_out0;
wire v$S_1569_out0;
wire v$S_1570_out0;
wire v$S_1571_out0;
wire v$S_1572_out0;
wire v$S_1573_out0;
wire v$S_1574_out0;
wire v$S_1575_out0;
wire v$S_1576_out0;
wire v$S_1577_out0;
wire v$S_1578_out0;
wire v$S_1579_out0;
wire v$S_1580_out0;
wire v$S_1581_out0;
wire v$S_1582_out0;
wire v$S_1583_out0;
wire v$S_1584_out0;
wire v$S_1585_out0;
wire v$S_1586_out0;
wire v$S_1587_out0;
wire v$S_1588_out0;
wire v$S_1589_out0;
wire v$S_1590_out0;
wire v$S_1591_out0;
wire v$S_1592_out0;
wire v$S_1593_out0;
wire v$S_1594_out0;
wire v$S_1595_out0;
wire v$S_1596_out0;
wire v$S_1597_out0;
wire v$S_1598_out0;
wire v$S_1599_out0;
wire v$S_1600_out0;
wire v$S_1601_out0;
wire v$S_1602_out0;
wire v$S_1603_out0;
wire v$S_1604_out0;
wire v$S_1605_out0;
wire v$S_1606_out0;
wire v$S_1607_out0;
wire v$S_1608_out0;
wire v$S_1609_out0;
wire v$S_1610_out0;
wire v$S_1611_out0;
wire v$S_1612_out0;
wire v$S_1613_out0;
wire v$S_1614_out0;
wire v$S_1615_out0;
wire v$S_1616_out0;
wire v$S_1617_out0;
wire v$S_1618_out0;
wire v$S_1619_out0;
wire v$S_1620_out0;
wire v$S_1621_out0;
wire v$S_1622_out0;
wire v$S_1623_out0;
wire v$S_1624_out0;
wire v$S_1625_out0;
wire v$S_1626_out0;
wire v$S_1627_out0;
wire v$S_1628_out0;
wire v$S_1629_out0;
wire v$S_1630_out0;
wire v$S_1631_out0;
wire v$S_1632_out0;
wire v$S_1633_out0;
wire v$S_1634_out0;
wire v$S_1635_out0;
wire v$S_1636_out0;
wire v$S_1637_out0;
wire v$S_1638_out0;
wire v$S_1639_out0;
wire v$S_1640_out0;
wire v$S_1641_out0;
wire v$S_1642_out0;
wire v$S_1643_out0;
wire v$S_1644_out0;
wire v$S_1645_out0;
wire v$S_1646_out0;
wire v$S_1647_out0;
wire v$S_1648_out0;
wire v$S_1649_out0;
wire v$S_1650_out0;
wire v$S_1651_out0;
wire v$S_1652_out0;
wire v$S_1653_out0;
wire v$S_1654_out0;
wire v$S_1655_out0;
wire v$S_1656_out0;
wire v$S_1657_out0;
wire v$S_1658_out0;
wire v$S_1659_out0;
wire v$S_1660_out0;
wire v$S_1661_out0;
wire v$S_1662_out0;
wire v$S_1663_out0;
wire v$S_1664_out0;
wire v$S_1665_out0;
wire v$S_1666_out0;
wire v$S_4665_out0;
wire v$S_4666_out0;
wire v$S_4667_out0;
wire v$S_4668_out0;
wire v$S_4669_out0;
wire v$S_4670_out0;
wire v$S_4671_out0;
wire v$S_4672_out0;
wire v$S_4673_out0;
wire v$S_4674_out0;
wire v$S_4675_out0;
wire v$S_4676_out0;
wire v$S_4677_out0;
wire v$S_4678_out0;
wire v$S_4679_out0;
wire v$S_4680_out0;
wire v$S_4681_out0;
wire v$S_4682_out0;
wire v$S_4683_out0;
wire v$S_4684_out0;
wire v$S_4685_out0;
wire v$S_4686_out0;
wire v$S_4687_out0;
wire v$S_4688_out0;
wire v$S_4689_out0;
wire v$S_4690_out0;
wire v$S_4691_out0;
wire v$S_4692_out0;
wire v$S_4693_out0;
wire v$S_4694_out0;
wire v$S_8863_out0;
wire v$S_8864_out0;
wire v$S_8865_out0;
wire v$S_8866_out0;
wire v$S_8867_out0;
wire v$S_8868_out0;
wire v$S_8869_out0;
wire v$S_8870_out0;
wire v$S_8871_out0;
wire v$S_8872_out0;
wire v$S_8873_out0;
wire v$S_8874_out0;
wire v$S_8875_out0;
wire v$S_8876_out0;
wire v$S_8877_out0;
wire v$S_8878_out0;
wire v$S_8879_out0;
wire v$S_8880_out0;
wire v$S_8881_out0;
wire v$S_8882_out0;
wire v$S_8883_out0;
wire v$S_8884_out0;
wire v$S_8885_out0;
wire v$S_8886_out0;
wire v$S_8887_out0;
wire v$S_8888_out0;
wire v$S_8889_out0;
wire v$S_8890_out0;
wire v$S_8891_out0;
wire v$S_8892_out0;
wire v$S_8893_out0;
wire v$S_8894_out0;
wire v$S_8895_out0;
wire v$S_8896_out0;
wire v$S_8897_out0;
wire v$S_8898_out0;
wire v$S_8899_out0;
wire v$S_8900_out0;
wire v$S_8901_out0;
wire v$S_8902_out0;
wire v$S_8903_out0;
wire v$S_8904_out0;
wire v$S_8905_out0;
wire v$S_8906_out0;
wire v$S_8907_out0;
wire v$S_8908_out0;
wire v$S_8909_out0;
wire v$S_8910_out0;
wire v$S_8911_out0;
wire v$S_8912_out0;
wire v$S_8913_out0;
wire v$S_8914_out0;
wire v$S_8915_out0;
wire v$S_8916_out0;
wire v$S_8917_out0;
wire v$S_8918_out0;
wire v$S_8919_out0;
wire v$S_8920_out0;
wire v$S_8921_out0;
wire v$S_8922_out0;
wire v$S_8923_out0;
wire v$S_8924_out0;
wire v$S_8925_out0;
wire v$S_8926_out0;
wire v$S_8927_out0;
wire v$S_8928_out0;
wire v$S_8929_out0;
wire v$S_8930_out0;
wire v$S_8931_out0;
wire v$S_8932_out0;
wire v$S_8933_out0;
wire v$S_8934_out0;
wire v$S_8935_out0;
wire v$S_8936_out0;
wire v$S_8937_out0;
wire v$S_8938_out0;
wire v$S_8939_out0;
wire v$S_8940_out0;
wire v$S_8941_out0;
wire v$S_8942_out0;
wire v$S_8943_out0;
wire v$S_8944_out0;
wire v$S_8945_out0;
wire v$S_8946_out0;
wire v$S_8947_out0;
wire v$S_8948_out0;
wire v$S_8949_out0;
wire v$S_8950_out0;
wire v$S_8951_out0;
wire v$S_8952_out0;
wire v$S_8953_out0;
wire v$S_8954_out0;
wire v$S_8955_out0;
wire v$S_8956_out0;
wire v$S_8957_out0;
wire v$S_8958_out0;
wire v$S_8959_out0;
wire v$S_8960_out0;
wire v$S_8961_out0;
wire v$S_8962_out0;
wire v$S_8963_out0;
wire v$S_8964_out0;
wire v$S_8965_out0;
wire v$S_8966_out0;
wire v$S_8967_out0;
wire v$S_8968_out0;
wire v$S_8969_out0;
wire v$S_8970_out0;
wire v$S_8971_out0;
wire v$S_8972_out0;
wire v$S_8973_out0;
wire v$S_8974_out0;
wire v$S_8975_out0;
wire v$S_8976_out0;
wire v$S_8977_out0;
wire v$S_8978_out0;
wire v$S_8979_out0;
wire v$S_8980_out0;
wire v$S_8981_out0;
wire v$S_8982_out0;
wire v$S_8983_out0;
wire v$S_8984_out0;
wire v$S_8985_out0;
wire v$S_8986_out0;
wire v$S_8987_out0;
wire v$S_8988_out0;
wire v$S_8989_out0;
wire v$S_8990_out0;
wire v$S_8991_out0;
wire v$S_8992_out0;
wire v$S_8993_out0;
wire v$S_8994_out0;
wire v$S_8995_out0;
wire v$S_8996_out0;
wire v$S_8997_out0;
wire v$S_8998_out0;
wire v$S_8999_out0;
wire v$S_9000_out0;
wire v$S_9001_out0;
wire v$S_9002_out0;
wire v$S_9003_out0;
wire v$S_9004_out0;
wire v$S_9005_out0;
wire v$S_9006_out0;
wire v$S_9007_out0;
wire v$S_9008_out0;
wire v$S_9009_out0;
wire v$S_9010_out0;
wire v$S_9011_out0;
wire v$S_9012_out0;
wire v$S_9013_out0;
wire v$S_9014_out0;
wire v$S_9015_out0;
wire v$S_9016_out0;
wire v$S_9017_out0;
wire v$S_9018_out0;
wire v$S_9019_out0;
wire v$S_9020_out0;
wire v$S_9021_out0;
wire v$S_9022_out0;
wire v$S_9023_out0;
wire v$S_9024_out0;
wire v$S_9025_out0;
wire v$S_9026_out0;
wire v$S_9027_out0;
wire v$S_9028_out0;
wire v$S_9029_out0;
wire v$S_9030_out0;
wire v$S_9031_out0;
wire v$S_9032_out0;
wire v$S_9033_out0;
wire v$S_9034_out0;
wire v$S_9035_out0;
wire v$S_9036_out0;
wire v$S_9037_out0;
wire v$S_9038_out0;
wire v$S_9039_out0;
wire v$S_9040_out0;
wire v$S_9041_out0;
wire v$S_9042_out0;
wire v$S_9043_out0;
wire v$S_9044_out0;
wire v$S_9045_out0;
wire v$S_9046_out0;
wire v$S_9047_out0;
wire v$S_9048_out0;
wire v$S_9049_out0;
wire v$S_9050_out0;
wire v$S_9051_out0;
wire v$S_9052_out0;
wire v$S_9053_out0;
wire v$S_9054_out0;
wire v$S_9055_out0;
wire v$S_9056_out0;
wire v$S_9057_out0;
wire v$S_9058_out0;
wire v$S_9059_out0;
wire v$S_9060_out0;
wire v$S_9061_out0;
wire v$S_9062_out0;
wire v$S_9063_out0;
wire v$S_9064_out0;
wire v$S_9065_out0;
wire v$S_9066_out0;
wire v$S_9067_out0;
wire v$S_9068_out0;
wire v$S_9069_out0;
wire v$S_9070_out0;
wire v$S_9071_out0;
wire v$S_9072_out0;
wire v$S_9073_out0;
wire v$S_9074_out0;
wire v$S_9075_out0;
wire v$S_9076_out0;
wire v$S_9077_out0;
wire v$S_9078_out0;
wire v$S_9079_out0;
wire v$S_9080_out0;
wire v$S_9081_out0;
wire v$S_9082_out0;
wire v$S_9083_out0;
wire v$S_9084_out0;
wire v$S_9085_out0;
wire v$S_9086_out0;
wire v$S_9087_out0;
wire v$S_9088_out0;
wire v$S_9089_out0;
wire v$S_9090_out0;
wire v$S_9091_out0;
wire v$S_9092_out0;
wire v$S_9093_out0;
wire v$S_9094_out0;
wire v$S_9095_out0;
wire v$S_9096_out0;
wire v$S_9097_out0;
wire v$S_9098_out0;
wire v$S_9099_out0;
wire v$S_9100_out0;
wire v$S_9101_out0;
wire v$S_9102_out0;
wire v$S_9103_out0;
wire v$S_9104_out0;
wire v$S_9105_out0;
wire v$S_9106_out0;
wire v$S_9107_out0;
wire v$S_9108_out0;
wire v$S_9109_out0;
wire v$S_9110_out0;
wire v$S_9111_out0;
wire v$S_9112_out0;
wire v$S_9113_out0;
wire v$S_9114_out0;
wire v$S_9115_out0;
wire v$S_9116_out0;
wire v$S_9117_out0;
wire v$S_9118_out0;
wire v$S_9119_out0;
wire v$S_9120_out0;
wire v$S_9121_out0;
wire v$S_9122_out0;
wire v$S_9123_out0;
wire v$S_9124_out0;
wire v$S_9125_out0;
wire v$S_9126_out0;
wire v$S_9127_out0;
wire v$S_9128_out0;
wire v$S_9129_out0;
wire v$S_9130_out0;
wire v$S_9131_out0;
wire v$S_9132_out0;
wire v$S_9133_out0;
wire v$S_9134_out0;
wire v$S_9135_out0;
wire v$S_9136_out0;
wire v$S_9137_out0;
wire v$S_9138_out0;
wire v$S_9139_out0;
wire v$S_9140_out0;
wire v$S_9141_out0;
wire v$S_9142_out0;
wire v$S_9143_out0;
wire v$S_9144_out0;
wire v$S_9145_out0;
wire v$S_9146_out0;
wire v$S_9147_out0;
wire v$S_9148_out0;
wire v$S_9149_out0;
wire v$S_9150_out0;
wire v$S_9151_out0;
wire v$S_9152_out0;
wire v$S_9153_out0;
wire v$S_9154_out0;
wire v$S_9155_out0;
wire v$S_9156_out0;
wire v$S_9157_out0;
wire v$S_9158_out0;
wire v$S_9159_out0;
wire v$S_9160_out0;
wire v$S_9161_out0;
wire v$S_9162_out0;
wire v$S_9163_out0;
wire v$S_9164_out0;
wire v$S_9165_out0;
wire v$S_9166_out0;
wire v$S_9167_out0;
wire v$S_9168_out0;
wire v$S_9169_out0;
wire v$S_9170_out0;
wire v$S_9171_out0;
wire v$S_9172_out0;
wire v$S_9173_out0;
wire v$S_9174_out0;
wire v$S_9175_out0;
wire v$S_9176_out0;
wire v$S_9177_out0;
wire v$S_9178_out0;
wire v$S_9179_out0;
wire v$S_9180_out0;
wire v$S_9181_out0;
wire v$S_9182_out0;
wire v$S_9183_out0;
wire v$S_9184_out0;
wire v$S_9185_out0;
wire v$S_9186_out0;
wire v$S_9187_out0;
wire v$S_9188_out0;
wire v$S_9189_out0;
wire v$S_9190_out0;
wire v$S_9191_out0;
wire v$S_9192_out0;
wire v$S_9193_out0;
wire v$S_9194_out0;
wire v$S_9195_out0;
wire v$S_9196_out0;
wire v$S_9197_out0;
wire v$S_9198_out0;
wire v$S_9199_out0;
wire v$S_9200_out0;
wire v$S_9201_out0;
wire v$S_9202_out0;
wire v$S_9203_out0;
wire v$S_9204_out0;
wire v$S_9205_out0;
wire v$S_9206_out0;
wire v$S_9207_out0;
wire v$S_9208_out0;
wire v$S_9209_out0;
wire v$S_9210_out0;
wire v$S_9211_out0;
wire v$S_9212_out0;
wire v$S_9213_out0;
wire v$S_9214_out0;
wire v$S_9215_out0;
wire v$S_9216_out0;
wire v$S_9217_out0;
wire v$S_9218_out0;
wire v$S_9219_out0;
wire v$S_9220_out0;
wire v$S_9221_out0;
wire v$S_9222_out0;
wire v$S_9223_out0;
wire v$S_9224_out0;
wire v$S_9225_out0;
wire v$S_9226_out0;
wire v$S_9227_out0;
wire v$S_9228_out0;
wire v$S_9229_out0;
wire v$S_9230_out0;
wire v$S_9231_out0;
wire v$S_9232_out0;
wire v$S_9233_out0;
wire v$S_9234_out0;
wire v$S_9235_out0;
wire v$S_9236_out0;
wire v$S_9237_out0;
wire v$S_9238_out0;
wire v$S_9239_out0;
wire v$S_9240_out0;
wire v$S_9241_out0;
wire v$S_9242_out0;
wire v$S_9243_out0;
wire v$S_9244_out0;
wire v$S_9245_out0;
wire v$S_9246_out0;
wire v$S_9247_out0;
wire v$S_9248_out0;
wire v$S_9249_out0;
wire v$S_9250_out0;
wire v$S_9251_out0;
wire v$S_9252_out0;
wire v$S_9253_out0;
wire v$S_9254_out0;
wire v$S_9255_out0;
wire v$S_9256_out0;
wire v$S_9257_out0;
wire v$S_9258_out0;
wire v$S_9259_out0;
wire v$S_9260_out0;
wire v$S_9261_out0;
wire v$S_9262_out0;
wire v$S_9263_out0;
wire v$S_9264_out0;
wire v$S_9265_out0;
wire v$S_9266_out0;
wire v$S_9267_out0;
wire v$S_9268_out0;
wire v$S_9269_out0;
wire v$S_9270_out0;
wire v$S_9271_out0;
wire v$S_9272_out0;
wire v$S_9273_out0;
wire v$S_9274_out0;
wire v$S_9275_out0;
wire v$S_9276_out0;
wire v$S_9277_out0;
wire v$S_9278_out0;
wire v$S_9279_out0;
wire v$S_9280_out0;
wire v$S_9281_out0;
wire v$S_9282_out0;
wire v$S_9283_out0;
wire v$S_9284_out0;
wire v$S_9285_out0;
wire v$S_9286_out0;
wire v$S_9287_out0;
wire v$S_9288_out0;
wire v$S_9289_out0;
wire v$S_9290_out0;
wire v$S_9291_out0;
wire v$S_9292_out0;
wire v$S_9293_out0;
wire v$S_9294_out0;
wire v$S_9295_out0;
wire v$S_9296_out0;
wire v$S_9297_out0;
wire v$S_9298_out0;
wire v$S_9299_out0;
wire v$S_9300_out0;
wire v$S_9301_out0;
wire v$S_9302_out0;
wire v$S_9303_out0;
wire v$S_9304_out0;
wire v$S_9305_out0;
wire v$S_9306_out0;
wire v$S_9307_out0;
wire v$S_9308_out0;
wire v$S_9309_out0;
wire v$S_9310_out0;
wire v$S_9311_out0;
wire v$S_9312_out0;
wire v$S_9313_out0;
wire v$S_9314_out0;
wire v$S_9315_out0;
wire v$S_9316_out0;
wire v$S_9317_out0;
wire v$S_9318_out0;
wire v$S_9319_out0;
wire v$S_9320_out0;
wire v$S_9321_out0;
wire v$S_9322_out0;
wire v$S_9323_out0;
wire v$S_9324_out0;
wire v$S_9325_out0;
wire v$S_9326_out0;
wire v$S_9327_out0;
wire v$S_9328_out0;
wire v$S_9329_out0;
wire v$S_9330_out0;
wire v$S_9331_out0;
wire v$S_9332_out0;
wire v$S_9333_out0;
wire v$S_9334_out0;
wire v$S_9335_out0;
wire v$S_9336_out0;
wire v$S_9337_out0;
wire v$S_9338_out0;
wire v$S_9339_out0;
wire v$S_9340_out0;
wire v$S_9341_out0;
wire v$S_9342_out0;
wire v$S_9343_out0;
wire v$S_9344_out0;
wire v$S_9345_out0;
wire v$S_9346_out0;
wire v$S_9347_out0;
wire v$S_9348_out0;
wire v$S_9349_out0;
wire v$S_9350_out0;
wire v$S_9351_out0;
wire v$S_9352_out0;
wire v$S_9353_out0;
wire v$S_9354_out0;
wire v$S_9355_out0;
wire v$S_9356_out0;
wire v$S_9357_out0;
wire v$S_9358_out0;
wire v$S_9359_out0;
wire v$S_9360_out0;
wire v$S_9361_out0;
wire v$S_9362_out0;
wire v$S_9363_out0;
wire v$S_9364_out0;
wire v$S_9365_out0;
wire v$S_9366_out0;
wire v$S_9367_out0;
wire v$S_9368_out0;
wire v$S_9369_out0;
wire v$S_9370_out0;
wire v$S_9371_out0;
wire v$S_9372_out0;
wire v$S_9373_out0;
wire v$S_9374_out0;
wire v$S_9375_out0;
wire v$S_9376_out0;
wire v$S_9377_out0;
wire v$S_9378_out0;
wire v$S_9379_out0;
wire v$S_9380_out0;
wire v$S_9381_out0;
wire v$S_9382_out0;
wire v$S_9383_out0;
wire v$S_9384_out0;
wire v$S_9385_out0;
wire v$S_9386_out0;
wire v$S_9387_out0;
wire v$S_9388_out0;
wire v$S_9389_out0;
wire v$S_9390_out0;
wire v$S_9391_out0;
wire v$S_9392_out0;
wire v$S_9393_out0;
wire v$S_9394_out0;
wire v$S_9395_out0;
wire v$S_9396_out0;
wire v$S_9397_out0;
wire v$S_9398_out0;
wire v$S_9399_out0;
wire v$S_9400_out0;
wire v$S_9401_out0;
wire v$S_9402_out0;
wire v$S_9403_out0;
wire v$S_9404_out0;
wire v$S_9405_out0;
wire v$S_9406_out0;
wire v$S_9407_out0;
wire v$S_9408_out0;
wire v$S_9409_out0;
wire v$S_9410_out0;
wire v$S_9411_out0;
wire v$S_9412_out0;
wire v$S_9413_out0;
wire v$S_9414_out0;
wire v$S_9415_out0;
wire v$S_9416_out0;
wire v$S_9417_out0;
wire v$S_9418_out0;
wire v$S_9419_out0;
wire v$S_9420_out0;
wire v$S_9421_out0;
wire v$S_9422_out0;
wire v$S_9423_out0;
wire v$S_9424_out0;
wire v$S_9425_out0;
wire v$S_9426_out0;
wire v$S_9427_out0;
wire v$S_9428_out0;
wire v$S_9429_out0;
wire v$S_9430_out0;
wire v$S_9431_out0;
wire v$S_9432_out0;
wire v$S_9433_out0;
wire v$S_9434_out0;
wire v$S_9435_out0;
wire v$S_9436_out0;
wire v$S_9437_out0;
wire v$S_9438_out0;
wire v$S_9439_out0;
wire v$S_9440_out0;
wire v$S_9441_out0;
wire v$S_9442_out0;
wire v$S_9443_out0;
wire v$S_9444_out0;
wire v$S_9445_out0;
wire v$S_9446_out0;
wire v$S_9447_out0;
wire v$S_9448_out0;
wire v$S_9449_out0;
wire v$S_9450_out0;
wire v$S_9451_out0;
wire v$S_9452_out0;
wire v$S_9453_out0;
wire v$S_9454_out0;
wire v$S_9455_out0;
wire v$S_9456_out0;
wire v$S_9457_out0;
wire v$S_9458_out0;
wire v$S_9459_out0;
wire v$S_9460_out0;
wire v$S_9461_out0;
wire v$S_9462_out0;
wire v$S_9463_out0;
wire v$S_9464_out0;
wire v$S_9465_out0;
wire v$S_9466_out0;
wire v$S_9467_out0;
wire v$S_9468_out0;
wire v$S_9469_out0;
wire v$S_9470_out0;
wire v$S_9471_out0;
wire v$S_9472_out0;
wire v$S_9473_out0;
wire v$S_9474_out0;
wire v$S_9475_out0;
wire v$S_9476_out0;
wire v$S_9477_out0;
wire v$S_9478_out0;
wire v$S_9479_out0;
wire v$S_9480_out0;
wire v$S_9481_out0;
wire v$S_9482_out0;
wire v$S_9483_out0;
wire v$S_9484_out0;
wire v$S_9485_out0;
wire v$S_9486_out0;
wire v$S_9487_out0;
wire v$S_9488_out0;
wire v$S_9489_out0;
wire v$S_9490_out0;
wire v$S_9491_out0;
wire v$S_9492_out0;
wire v$S_9493_out0;
wire v$S_9494_out0;
wire v$S_9495_out0;
wire v$S_9496_out0;
wire v$S_9497_out0;
wire v$S_9498_out0;
wire v$S_9499_out0;
wire v$S_9500_out0;
wire v$S_9501_out0;
wire v$S_9502_out0;
wire v$S_9503_out0;
wire v$S_9504_out0;
wire v$S_9505_out0;
wire v$S_9506_out0;
wire v$S_9507_out0;
wire v$S_9508_out0;
wire v$S_9509_out0;
wire v$S_9510_out0;
wire v$S_9511_out0;
wire v$S_9512_out0;
wire v$S_9513_out0;
wire v$S_9514_out0;
wire v$S_9515_out0;
wire v$S_9516_out0;
wire v$S_9517_out0;
wire v$S_9518_out0;
wire v$S_9519_out0;
wire v$S_9520_out0;
wire v$S_9521_out0;
wire v$S_9522_out0;
wire v$S_9523_out0;
wire v$S_9524_out0;
wire v$S_9525_out0;
wire v$S_9526_out0;
wire v$S_9527_out0;
wire v$S_9528_out0;
wire v$S_9529_out0;
wire v$S_9530_out0;
wire v$S_9531_out0;
wire v$S_9532_out0;
wire v$S_9533_out0;
wire v$S_9534_out0;
wire v$S_9535_out0;
wire v$S_9536_out0;
wire v$S_9537_out0;
wire v$S_9538_out0;
wire v$S_9539_out0;
wire v$S_9540_out0;
wire v$S_9541_out0;
wire v$S_9542_out0;
wire v$S_9543_out0;
wire v$S_9544_out0;
wire v$S_9545_out0;
wire v$S_9546_out0;
wire v$S_9547_out0;
wire v$S_9548_out0;
wire v$S_9549_out0;
wire v$S_9550_out0;
wire v$S_9551_out0;
wire v$S_9552_out0;
wire v$S_9553_out0;
wire v$S_9554_out0;
wire v$S_9555_out0;
wire v$S_9556_out0;
wire v$S_9557_out0;
wire v$S_9558_out0;
wire v$S_9559_out0;
wire v$S_9560_out0;
wire v$S_9561_out0;
wire v$S_9562_out0;
wire v$S_9563_out0;
wire v$S_9564_out0;
wire v$S_9565_out0;
wire v$S_9566_out0;
wire v$S_9567_out0;
wire v$S_9568_out0;
wire v$S_9569_out0;
wire v$S_9570_out0;
wire v$S_9571_out0;
wire v$S_9572_out0;
wire v$S_9573_out0;
wire v$S_9574_out0;
wire v$S_9575_out0;
wire v$S_9576_out0;
wire v$S_9577_out0;
wire v$S_9578_out0;
wire v$S_9579_out0;
wire v$S_9580_out0;
wire v$S_9581_out0;
wire v$S_9582_out0;
wire v$S_9583_out0;
wire v$S_9584_out0;
wire v$S_9585_out0;
wire v$S_9586_out0;
wire v$S_9587_out0;
wire v$S_9588_out0;
wire v$S_9589_out0;
wire v$S_9590_out0;
wire v$S_9591_out0;
wire v$S_9592_out0;
wire v$S_9593_out0;
wire v$S_9594_out0;
wire v$S_9595_out0;
wire v$S_9596_out0;
wire v$S_9597_out0;
wire v$S_9598_out0;
wire v$S_9599_out0;
wire v$S_9600_out0;
wire v$S_9601_out0;
wire v$S_9602_out0;
wire v$S_9603_out0;
wire v$S_9604_out0;
wire v$S_9605_out0;
wire v$S_9606_out0;
wire v$S_9607_out0;
wire v$S_9608_out0;
wire v$S_9609_out0;
wire v$S_9610_out0;
wire v$S_9611_out0;
wire v$S_9612_out0;
wire v$S_9613_out0;
wire v$S_9614_out0;
wire v$S_9615_out0;
wire v$S_9616_out0;
wire v$S_9617_out0;
wire v$S_9618_out0;
wire v$S_9619_out0;
wire v$S_9620_out0;
wire v$S_9621_out0;
wire v$S_9622_out0;
wire v$S_9623_out0;
wire v$S_9624_out0;
wire v$S_9625_out0;
wire v$S_9626_out0;
wire v$S_9627_out0;
wire v$S_9628_out0;
wire v$S_9629_out0;
wire v$S_9630_out0;
wire v$S_9631_out0;
wire v$S_9632_out0;
wire v$S_9633_out0;
wire v$S_9634_out0;
wire v$S_9635_out0;
wire v$S_9636_out0;
wire v$S_9637_out0;
wire v$S_9638_out0;
wire v$S_9639_out0;
wire v$S_9640_out0;
wire v$S_9641_out0;
wire v$S_9642_out0;
wire v$S_9643_out0;
wire v$S_9644_out0;
wire v$S_9645_out0;
wire v$S_9646_out0;
wire v$S_9647_out0;
wire v$S_9648_out0;
wire v$S_9649_out0;
wire v$S_9650_out0;
wire v$S_9651_out0;
wire v$S_9652_out0;
wire v$S_9653_out0;
wire v$S_9654_out0;
wire v$S_9655_out0;
wire v$S_9656_out0;
wire v$S_9657_out0;
wire v$S_9658_out0;
wire v$S_9659_out0;
wire v$S_9660_out0;
wire v$S_9661_out0;
wire v$S_9662_out0;
wire v$S_9663_out0;
wire v$S_9664_out0;
wire v$S_9665_out0;
wire v$S_9666_out0;
wire v$S_9667_out0;
wire v$S_9668_out0;
wire v$S_9669_out0;
wire v$S_9670_out0;
wire v$S_9671_out0;
wire v$S_9672_out0;
wire v$S_9673_out0;
wire v$S_9674_out0;
wire v$S_9675_out0;
wire v$S_9676_out0;
wire v$S_9677_out0;
wire v$S_9678_out0;
wire v$S_9679_out0;
wire v$S_9680_out0;
wire v$S_9681_out0;
wire v$S_9682_out0;
wire v$S_9683_out0;
wire v$S_9684_out0;
wire v$S_9685_out0;
wire v$S_9686_out0;
wire v$S_9687_out0;
wire v$S_9688_out0;
wire v$S_9689_out0;
wire v$S_9690_out0;
wire v$S_9691_out0;
wire v$S_9692_out0;
wire v$S_9693_out0;
wire v$S_9694_out0;
wire v$S_9695_out0;
wire v$S_9696_out0;
wire v$S_9697_out0;
wire v$S_9698_out0;
wire v$S_9699_out0;
wire v$S_9700_out0;
wire v$S_9701_out0;
wire v$S_9702_out0;
wire v$S_9703_out0;
wire v$S_9704_out0;
wire v$S_9705_out0;
wire v$S_9706_out0;
wire v$S_9707_out0;
wire v$S_9708_out0;
wire v$S_9709_out0;
wire v$S_9710_out0;
wire v$S_9711_out0;
wire v$S_9712_out0;
wire v$S_9713_out0;
wire v$S_9714_out0;
wire v$S_9715_out0;
wire v$S_9716_out0;
wire v$S_9717_out0;
wire v$S_9718_out0;
wire v$S_9719_out0;
wire v$S_9720_out0;
wire v$S_9721_out0;
wire v$S_9722_out0;
wire v$S_9723_out0;
wire v$S_9724_out0;
wire v$S_9725_out0;
wire v$S_9726_out0;
wire v$S_9727_out0;
wire v$S_9728_out0;
wire v$S_9729_out0;
wire v$S_9730_out0;
wire v$S_9731_out0;
wire v$S_9732_out0;
wire v$S_9733_out0;
wire v$S_9734_out0;
wire v$S_9735_out0;
wire v$S_9736_out0;
wire v$S_9737_out0;
wire v$S_9738_out0;
wire v$S_9739_out0;
wire v$S_9740_out0;
wire v$S_9741_out0;
wire v$S_9742_out0;
wire v$S_9743_out0;
wire v$S_9744_out0;
wire v$S_9745_out0;
wire v$S_9746_out0;
wire v$S_9747_out0;
wire v$S_9748_out0;
wire v$S_9749_out0;
wire v$S_9750_out0;
wire v$S_9751_out0;
wire v$S_9752_out0;
wire v$S_9753_out0;
wire v$S_9754_out0;
wire v$S_9755_out0;
wire v$S_9756_out0;
wire v$S_9757_out0;
wire v$S_9758_out0;
wire v$S_9759_out0;
wire v$S_9760_out0;
wire v$S_9761_out0;
wire v$S_9762_out0;
wire v$S_9763_out0;
wire v$S_9764_out0;
wire v$S_9765_out0;
wire v$S_9766_out0;
wire v$S_9767_out0;
wire v$S_9768_out0;
wire v$S_9769_out0;
wire v$S_9770_out0;
wire v$S_9771_out0;
wire v$S_9772_out0;
wire v$S_9773_out0;
wire v$S_9774_out0;
wire v$S_9775_out0;
wire v$S_9776_out0;
wire v$S_9777_out0;
wire v$S_9778_out0;
wire v$S_9779_out0;
wire v$S_9780_out0;
wire v$S_9781_out0;
wire v$S_9782_out0;
wire v$S_9783_out0;
wire v$S_9784_out0;
wire v$S_9785_out0;
wire v$S_9786_out0;
wire v$S_9787_out0;
wire v$S_9788_out0;
wire v$S_9789_out0;
wire v$S_9790_out0;
wire v$TRANSMIT$INSTRUCTION_1713_out0;
wire v$TST_3819_out0;
wire v$TST_3820_out0;
wire v$TST_409_out0;
wire v$TST_410_out0;
wire v$TST_8735_out0;
wire v$TST_8736_out0;
wire v$TX$IN$PROGRESS_13634_out0;
wire v$TX$IN$PROGRESS_235_out0;
wire v$TX$INSTRUCTION0_1762_out0;
wire v$TX$INSTRUCTION1_1169_out0;
wire v$TX$INSTRUCTION_10501_out0;
wire v$TX$INSTRUCTION_13631_out0;
wire v$TX$INSTRUCTION_13659_out0;
wire v$TX$INSTRUCTION_13660_out0;
wire v$TX$INSTRUCTION_2825_out0;
wire v$TX$INSTRUCTION_453_out0;
wire v$TX$INSTRUCTION_62_out0;
wire v$TX$INSTRUCTION_63_out0;
wire v$TX$INSTRUCTION_6875_out0;
wire v$TX$INSTRUCTION_7012_out0;
wire v$TX$INSTRUCTION_7013_out0;
wire v$TX$INSTUCTION0_228_out0;
wire v$TX$INSTUCTION1_4859_out0;
wire v$TX$INST_10827_out0;
wire v$TX$INST_10828_out0;
wire v$TX$INST_11239_out0;
wire v$TX$OVERFLOW_10481_out0;
wire v$TX$OVERFLOW_13294_out0;
wire v$TX$OVERFLOW_500_out0;
wire v$TX$PROGRESS_8645_out0;
wire v$TX$inst0_608_out0;
wire v$UART_10516_out0;
wire v$UART_10517_out0;
wire v$UART_10825_out0;
wire v$UART_10826_out0;
wire v$UART_11128_out0;
wire v$UART_11129_out0;
wire v$UART_1823_out0;
wire v$UART_1824_out0;
wire v$UART_3893_out0;
wire v$UART_3894_out0;
wire v$UNDERFLOW_6916_out0;
wire v$UNDERFLOW_6917_out0;
wire v$UNNOTUSED_11220_out0;
wire v$UNNOTUSED_11221_out0;
wire v$UNUSED1_3016_out0;
wire v$UNUSED1_3017_out0;
wire v$UNUSED1_3220_out0;
wire v$UNUSED2_2193_out0;
wire v$UNUSED2_2194_out0;
wire v$UNUSED2_2424_out0;
wire v$UNUSED3_1681_out0;
wire v$UNUSED_123_out0;
wire v$UNUSED_339_out0;
wire v$UNUSED_340_out0;
wire v$U_10469_out0;
wire v$U_10470_out0;
wire v$W$EN_6878_out0;
wire v$W$EN_6879_out0;
wire v$WEN$MULTI_10381_out0;
wire v$WEN$MULTI_10382_out0;
wire v$WEN$MULTI_2388_out0;
wire v$WEN$MULTI_2389_out0;
wire v$WEN$MULTI_35_out0;
wire v$WEN$MULTI_36_out0;
wire v$WEN$RAM_7079_out0;
wire v$WEN$RAM_7080_out0;
wire v$WEN0_13300_out0;
wire v$WEN0_2588_out0;
wire v$WEN0_2646_out0;
wire v$WEN1_7716_out0;
wire v$WEN1_8763_out0;
wire v$WEN3_1690_out0;
wire v$WEN3_1691_out0;
wire v$WENALU_10866_out0;
wire v$WENALU_10867_out0;
wire v$WENALU_8659_out0;
wire v$WENALU_8660_out0;
wire v$WENLDST_13755_out0;
wire v$WENLDST_13756_out0;
wire v$WENLDST_2682_out0;
wire v$WENLDST_2683_out0;
wire v$WENLS_11260_out0;
wire v$WENLS_11261_out0;
wire v$WENLS_600_out0;
wire v$WENLS_601_out0;
wire v$WENMULTI_11206_out0;
wire v$WENMULTI_11207_out0;
wire v$WENRAM_2326_out0;
wire v$WENRAM_2327_out0;
wire v$WENRAM_4650_out0;
wire v$WENRAM_4651_out0;
wire v$WEN_11038_out0;
wire v$WEN_11039_out0;
wire v$WEN_2154_out0;
wire v$WEN_2765_out0;
wire v$WEN_2766_out0;
wire v$WEN_3204_out0;
wire v$WRITE$EN_13653_out0;
wire v$WRITE$EN_13654_out0;
wire v$WWNELS0_385_out0;
wire v$WWNELS1_47_out0;
wire v$Wen1_10312_out0;
wire v$_0_out0;
wire v$_10377_out0;
wire v$_10378_out0;
wire v$_10379_out0;
wire v$_10380_out0;
wire v$_10385_out0;
wire v$_10386_out0;
wire v$_10387_out0;
wire v$_10388_out0;
wire v$_10409_out0;
wire v$_10410_out0;
wire v$_10411_out0;
wire v$_10412_out0;
wire v$_10413_out0;
wire v$_10414_out0;
wire v$_10415_out0;
wire v$_10416_out0;
wire v$_10417_out0;
wire v$_10418_out0;
wire v$_10419_out0;
wire v$_10420_out0;
wire v$_10421_out0;
wire v$_10422_out0;
wire v$_10423_out0;
wire v$_10424_out0;
wire v$_10425_out0;
wire v$_10426_out0;
wire v$_10427_out0;
wire v$_10428_out0;
wire v$_10429_out0;
wire v$_10430_out0;
wire v$_10431_out0;
wire v$_10432_out0;
wire v$_10433_out0;
wire v$_10434_out0;
wire v$_10435_out0;
wire v$_10436_out0;
wire v$_10437_out0;
wire v$_10438_out0;
wire v$_10472_out0;
wire v$_10473_out0;
wire v$_10479_out0;
wire v$_10480_out0;
wire v$_10490_out1;
wire v$_10491_out1;
wire v$_10536_out0;
wire v$_10537_out0;
wire v$_10538_out0;
wire v$_10539_out0;
wire v$_10695_out0;
wire v$_10696_out0;
wire v$_10697_out0;
wire v$_10698_out0;
wire v$_10717_out0;
wire v$_10718_out0;
wire v$_10719_out0;
wire v$_10720_out0;
wire v$_10721_out0;
wire v$_10722_out0;
wire v$_10723_out0;
wire v$_10724_out0;
wire v$_10725_out0;
wire v$_10726_out0;
wire v$_10727_out0;
wire v$_10728_out0;
wire v$_10729_out0;
wire v$_10730_out0;
wire v$_10731_out0;
wire v$_10732_out0;
wire v$_10733_out0;
wire v$_10734_out0;
wire v$_10735_out0;
wire v$_10736_out0;
wire v$_10737_out0;
wire v$_10738_out0;
wire v$_10739_out0;
wire v$_10740_out0;
wire v$_10741_out0;
wire v$_10742_out0;
wire v$_10743_out0;
wire v$_10744_out0;
wire v$_10745_out0;
wire v$_10746_out0;
wire v$_10747_out0;
wire v$_10748_out0;
wire v$_10777_out0;
wire v$_10778_out0;
wire v$_10779_out0;
wire v$_10780_out0;
wire v$_10785_out0;
wire v$_10786_out0;
wire v$_10808_out0;
wire v$_10809_out0;
wire v$_10823_out0;
wire v$_10824_out0;
wire v$_10862_out0;
wire v$_10863_out0;
wire v$_10864_out0;
wire v$_10865_out0;
wire v$_10868_out1;
wire v$_10869_out1;
wire v$_10874_out0;
wire v$_10875_out0;
wire v$_10876_out0;
wire v$_10877_out0;
wire v$_10878_out0;
wire v$_10879_out0;
wire v$_10880_out0;
wire v$_10881_out0;
wire v$_10882_out0;
wire v$_10883_out0;
wire v$_10884_out0;
wire v$_10885_out0;
wire v$_10886_out0;
wire v$_10887_out0;
wire v$_10888_out0;
wire v$_10889_out0;
wire v$_10890_out0;
wire v$_10891_out0;
wire v$_10892_out0;
wire v$_10893_out0;
wire v$_10894_out0;
wire v$_10895_out0;
wire v$_10896_out0;
wire v$_10897_out0;
wire v$_10898_out0;
wire v$_10899_out0;
wire v$_10900_out0;
wire v$_10901_out0;
wire v$_10902_out0;
wire v$_10903_out0;
wire v$_10910_out0;
wire v$_10911_out0;
wire v$_11001_out0;
wire v$_11002_out0;
wire v$_11003_out0;
wire v$_11004_out0;
wire v$_11005_out0;
wire v$_11006_out0;
wire v$_11007_out0;
wire v$_11008_out0;
wire v$_11009_out0;
wire v$_11010_out0;
wire v$_11011_out0;
wire v$_11012_out0;
wire v$_11013_out0;
wire v$_11014_out0;
wire v$_11015_out0;
wire v$_11016_out0;
wire v$_11017_out0;
wire v$_11018_out0;
wire v$_11019_out0;
wire v$_11020_out0;
wire v$_11021_out0;
wire v$_11022_out0;
wire v$_11023_out0;
wire v$_11024_out0;
wire v$_11025_out0;
wire v$_11026_out0;
wire v$_11027_out0;
wire v$_11028_out0;
wire v$_11029_out0;
wire v$_11030_out0;
wire v$_11098_out0;
wire v$_11099_out0;
wire v$_11100_out0;
wire v$_11101_out0;
wire v$_11102_out0;
wire v$_11103_out0;
wire v$_11104_out0;
wire v$_11105_out0;
wire v$_11106_out0;
wire v$_11107_out0;
wire v$_11108_out0;
wire v$_11109_out0;
wire v$_11110_out0;
wire v$_11111_out0;
wire v$_11112_out0;
wire v$_11113_out0;
wire v$_11114_out0;
wire v$_11115_out0;
wire v$_11116_out0;
wire v$_11117_out0;
wire v$_11118_out0;
wire v$_11119_out0;
wire v$_11120_out0;
wire v$_11121_out0;
wire v$_11122_out0;
wire v$_11123_out0;
wire v$_11124_out0;
wire v$_11125_out0;
wire v$_11126_out0;
wire v$_11127_out0;
wire v$_11149_out0;
wire v$_11150_out0;
wire v$_11151_out0;
wire v$_11152_out0;
wire v$_11212_out0;
wire v$_11213_out0;
wire v$_11242_out0;
wire v$_11243_out0;
wire v$_11294_out1;
wire v$_11295_out1;
wire v$_1176_out0;
wire v$_1177_out0;
wire v$_1193_out0;
wire v$_1194_out0;
wire v$_13251_out0;
wire v$_13252_out0;
wire v$_13384_out0;
wire v$_13385_out0;
wire v$_13386_out0;
wire v$_13387_out0;
wire v$_13392_out0;
wire v$_13393_out0;
wire v$_13396_out0;
wire v$_13397_out0;
wire v$_13399_out0;
wire v$_13400_out0;
wire v$_13401_out0;
wire v$_13402_out0;
wire v$_13403_out0;
wire v$_13404_out0;
wire v$_13405_out0;
wire v$_13406_out0;
wire v$_13407_out0;
wire v$_13408_out0;
wire v$_13409_out0;
wire v$_13410_out0;
wire v$_13411_out0;
wire v$_13412_out0;
wire v$_13413_out0;
wire v$_13414_out0;
wire v$_13415_out0;
wire v$_13416_out0;
wire v$_13417_out0;
wire v$_13418_out0;
wire v$_13419_out0;
wire v$_13420_out0;
wire v$_13421_out0;
wire v$_13422_out0;
wire v$_13423_out0;
wire v$_13424_out0;
wire v$_13425_out0;
wire v$_13426_out0;
wire v$_13427_out0;
wire v$_13428_out0;
wire v$_13435_out0;
wire v$_13436_out0;
wire v$_13448_out0;
wire v$_13449_out0;
wire v$_13450_out0;
wire v$_13451_out0;
wire v$_13452_out0;
wire v$_13453_out0;
wire v$_13454_out0;
wire v$_13455_out0;
wire v$_13456_out0;
wire v$_13457_out0;
wire v$_13458_out0;
wire v$_13459_out0;
wire v$_13460_out0;
wire v$_13461_out0;
wire v$_13462_out0;
wire v$_13463_out0;
wire v$_13464_out0;
wire v$_13465_out0;
wire v$_13466_out0;
wire v$_13467_out0;
wire v$_13468_out0;
wire v$_13469_out0;
wire v$_13470_out0;
wire v$_13471_out0;
wire v$_13472_out0;
wire v$_13473_out0;
wire v$_13474_out0;
wire v$_13475_out0;
wire v$_13476_out0;
wire v$_13477_out0;
wire v$_13512_out0;
wire v$_13513_out0;
wire v$_13514_out0;
wire v$_13515_out0;
wire v$_13552_out0;
wire v$_13553_out0;
wire v$_13554_out0;
wire v$_13555_out0;
wire v$_13562_out0;
wire v$_13563_out0;
wire v$_13601_out0;
wire v$_13602_out0;
wire v$_13627_out0;
wire v$_13628_out0;
wire v$_13629_out0;
wire v$_13630_out0;
wire v$_13715_out0;
wire v$_13716_out0;
wire v$_13717_out0;
wire v$_13718_out0;
wire v$_13719_out0;
wire v$_13720_out0;
wire v$_13721_out0;
wire v$_13722_out0;
wire v$_13723_out0;
wire v$_13724_out0;
wire v$_13725_out0;
wire v$_13726_out0;
wire v$_13727_out0;
wire v$_13728_out0;
wire v$_13729_out0;
wire v$_13730_out0;
wire v$_13731_out0;
wire v$_13732_out0;
wire v$_13733_out0;
wire v$_13734_out0;
wire v$_13735_out0;
wire v$_13736_out0;
wire v$_13737_out0;
wire v$_13738_out0;
wire v$_13739_out0;
wire v$_13740_out0;
wire v$_13741_out0;
wire v$_13742_out0;
wire v$_13743_out0;
wire v$_13744_out0;
wire v$_1692_out0;
wire v$_1693_out0;
wire v$_1694_out0;
wire v$_1695_out0;
wire v$_171_out0;
wire v$_1722_out0;
wire v$_1723_out0;
wire v$_1724_out0;
wire v$_1725_out0;
wire v$_1728_out0;
wire v$_1729_out0;
wire v$_172_out0;
wire v$_1747_out0;
wire v$_1748_out0;
wire v$_1749_out0;
wire v$_1750_out0;
wire v$_1773_out0;
wire v$_1774_out0;
wire v$_1775_out0;
wire v$_1776_out0;
wire v$_1777_out0;
wire v$_1778_out0;
wire v$_1779_out0;
wire v$_1780_out0;
wire v$_1781_out0;
wire v$_1782_out0;
wire v$_1783_out0;
wire v$_1784_out0;
wire v$_1785_out0;
wire v$_1786_out0;
wire v$_1787_out0;
wire v$_1788_out0;
wire v$_1789_out0;
wire v$_1790_out0;
wire v$_1791_out0;
wire v$_1792_out0;
wire v$_1793_out0;
wire v$_1794_out0;
wire v$_1795_out0;
wire v$_1796_out0;
wire v$_1797_out0;
wire v$_1798_out0;
wire v$_1799_out0;
wire v$_179_out0;
wire v$_1800_out0;
wire v$_1801_out0;
wire v$_1802_out0;
wire v$_180_out0;
wire v$_186_out0;
wire v$_1875_out0;
wire v$_1876_out0;
wire v$_187_out0;
wire v$_1893_out0;
wire v$_1894_out0;
wire v$_1895_out0;
wire v$_1896_out0;
wire v$_1904_out0;
wire v$_1905_out0;
wire v$_192_out0;
wire v$_193_out0;
wire v$_194_out0;
wire v$_195_out0;
wire v$_1975_out0;
wire v$_1976_out0;
wire v$_1977_out0;
wire v$_1978_out0;
wire v$_1979_out0;
wire v$_1980_out0;
wire v$_1981_out0;
wire v$_1982_out0;
wire v$_1983_out0;
wire v$_1984_out0;
wire v$_1985_out0;
wire v$_1986_out0;
wire v$_1987_out0;
wire v$_1988_out0;
wire v$_1989_out0;
wire v$_198_out0;
wire v$_1990_out0;
wire v$_1991_out0;
wire v$_1992_out0;
wire v$_1993_out0;
wire v$_1994_out0;
wire v$_1995_out0;
wire v$_1996_out0;
wire v$_1997_out0;
wire v$_1998_out0;
wire v$_1999_out0;
wire v$_199_out0;
wire v$_1_out0;
wire v$_2000_out0;
wire v$_2001_out0;
wire v$_2002_out0;
wire v$_2003_out0;
wire v$_2004_out0;
wire v$_2022_out0;
wire v$_2023_out0;
wire v$_2063_out0;
wire v$_2064_out0;
wire v$_2065_out0;
wire v$_2066_out0;
wire v$_2067_out0;
wire v$_2068_out0;
wire v$_2069_out0;
wire v$_2070_out0;
wire v$_2071_out0;
wire v$_2072_out0;
wire v$_2073_out0;
wire v$_2074_out0;
wire v$_2075_out0;
wire v$_2076_out0;
wire v$_2077_out0;
wire v$_2078_out0;
wire v$_2079_out0;
wire v$_2080_out0;
wire v$_2081_out0;
wire v$_2082_out0;
wire v$_2083_out0;
wire v$_2084_out0;
wire v$_2085_out0;
wire v$_2086_out0;
wire v$_2087_out0;
wire v$_2088_out0;
wire v$_2089_out0;
wire v$_2090_out0;
wire v$_2091_out0;
wire v$_2092_out0;
wire v$_2093_out0;
wire v$_2094_out0;
wire v$_2095_out0;
wire v$_2096_out0;
wire v$_2150_out0;
wire v$_2151_out0;
wire v$_2152_out0;
wire v$_2153_out0;
wire v$_2155_out0;
wire v$_2156_out0;
wire v$_2157_out0;
wire v$_2158_out0;
wire v$_2159_out0;
wire v$_2160_out0;
wire v$_2161_out0;
wire v$_2162_out0;
wire v$_2163_out0;
wire v$_2164_out0;
wire v$_2165_out0;
wire v$_2166_out0;
wire v$_2167_out0;
wire v$_2168_out0;
wire v$_2169_out0;
wire v$_2170_out0;
wire v$_2171_out0;
wire v$_2172_out0;
wire v$_2173_out0;
wire v$_2174_out0;
wire v$_2175_out0;
wire v$_2176_out0;
wire v$_2177_out0;
wire v$_2178_out0;
wire v$_2179_out0;
wire v$_2180_out0;
wire v$_2181_out0;
wire v$_2182_out0;
wire v$_2183_out0;
wire v$_2184_out0;
wire v$_2195_out0;
wire v$_2196_out0;
wire v$_2197_out0;
wire v$_2198_out0;
wire v$_2199_out0;
wire v$_2200_out0;
wire v$_2201_out0;
wire v$_2202_out0;
wire v$_2203_out0;
wire v$_2204_out0;
wire v$_2205_out0;
wire v$_2206_out0;
wire v$_2207_out0;
wire v$_2208_out0;
wire v$_2209_out0;
wire v$_2210_out0;
wire v$_2211_out0;
wire v$_2212_out0;
wire v$_2213_out0;
wire v$_2214_out0;
wire v$_2215_out0;
wire v$_2216_out0;
wire v$_2217_out0;
wire v$_2218_out0;
wire v$_2219_out0;
wire v$_2220_out0;
wire v$_2221_out0;
wire v$_2222_out0;
wire v$_2268_out0;
wire v$_2269_out0;
wire v$_2273_out0;
wire v$_2274_out0;
wire v$_2275_out0;
wire v$_2276_out0;
wire v$_2277_out0;
wire v$_2278_out0;
wire v$_2279_out0;
wire v$_2280_out0;
wire v$_2281_out0;
wire v$_2282_out0;
wire v$_2283_out0;
wire v$_2284_out0;
wire v$_2285_out0;
wire v$_2286_out0;
wire v$_2287_out0;
wire v$_2288_out0;
wire v$_2289_out0;
wire v$_2290_out0;
wire v$_2291_out0;
wire v$_2292_out0;
wire v$_2293_out0;
wire v$_2294_out0;
wire v$_2295_out0;
wire v$_2296_out0;
wire v$_2297_out0;
wire v$_2298_out0;
wire v$_2299_out0;
wire v$_2300_out0;
wire v$_2301_out0;
wire v$_2302_out0;
wire v$_2418_out0;
wire v$_2419_out0;
wire v$_2420_out0;
wire v$_2421_out0;
wire v$_2422_out0;
wire v$_2423_out0;
wire v$_2430_out0;
wire v$_2431_out0;
wire v$_2462_out0;
wire v$_2463_out0;
wire v$_2467_out0;
wire v$_2468_out0;
wire v$_2470_out0;
wire v$_2471_out0;
wire v$_2502_out0;
wire v$_2503_out0;
wire v$_2504_out0;
wire v$_2505_out0;
wire v$_2506_out0;
wire v$_2507_out0;
wire v$_2508_out0;
wire v$_2509_out0;
wire v$_2510_out0;
wire v$_2511_out0;
wire v$_2512_out0;
wire v$_2513_out0;
wire v$_2514_out0;
wire v$_2515_out0;
wire v$_2516_out0;
wire v$_2517_out0;
wire v$_2518_out0;
wire v$_2519_out0;
wire v$_2520_out0;
wire v$_2521_out0;
wire v$_2522_out0;
wire v$_2523_out0;
wire v$_2524_out0;
wire v$_2525_out0;
wire v$_2526_out0;
wire v$_2527_out0;
wire v$_2528_out0;
wire v$_2529_out0;
wire v$_2530_out0;
wire v$_2531_out0;
wire v$_2692_out0;
wire v$_2693_out0;
wire v$_2726_out0;
wire v$_2727_out0;
wire v$_2728_out0;
wire v$_2729_out0;
wire v$_2730_out0;
wire v$_2731_out0;
wire v$_2732_out0;
wire v$_2733_out0;
wire v$_2734_out0;
wire v$_2735_out0;
wire v$_2736_out0;
wire v$_2737_out0;
wire v$_2738_out0;
wire v$_2739_out0;
wire v$_2740_out0;
wire v$_2741_out0;
wire v$_2742_out0;
wire v$_2743_out0;
wire v$_2744_out0;
wire v$_2745_out0;
wire v$_2746_out0;
wire v$_2747_out0;
wire v$_2748_out0;
wire v$_2749_out0;
wire v$_2750_out0;
wire v$_2751_out0;
wire v$_2752_out0;
wire v$_2753_out0;
wire v$_2754_out0;
wire v$_2755_out0;
wire v$_2760_out0;
wire v$_2761_out0;
wire v$_2762_out0;
wire v$_2763_out0;
wire v$_2831_out0;
wire v$_2831_out1;
wire v$_2832_out0;
wire v$_2832_out1;
wire v$_2860_out0;
wire v$_2861_out0;
wire v$_2875_out0;
wire v$_2876_out0;
wire v$_2877_out0;
wire v$_2878_out0;
wire v$_2879_out0;
wire v$_287_out0;
wire v$_2880_out0;
wire v$_2881_out0;
wire v$_2882_out0;
wire v$_2889_out0;
wire v$_288_out0;
wire v$_2890_out0;
wire v$_2943_out0;
wire v$_2944_out0;
wire v$_2959_out0;
wire v$_2973_out0;
wire v$_2974_out0;
wire v$_2983_out0;
wire v$_2983_out1;
wire v$_2984_out0;
wire v$_2985_out0;
wire v$_2986_out0;
wire v$_2987_out0;
wire v$_2988_out0;
wire v$_2989_out0;
wire v$_2990_out0;
wire v$_2991_out0;
wire v$_2992_out0;
wire v$_2993_out0;
wire v$_2994_out0;
wire v$_2995_out0;
wire v$_2996_out0;
wire v$_2997_out0;
wire v$_2998_out0;
wire v$_2999_out0;
wire v$_2_out0;
wire v$_3000_out0;
wire v$_3001_out0;
wire v$_3002_out0;
wire v$_3003_out0;
wire v$_3004_out0;
wire v$_3005_out0;
wire v$_3006_out0;
wire v$_3007_out0;
wire v$_3008_out0;
wire v$_3009_out0;
wire v$_3010_out0;
wire v$_3011_out0;
wire v$_3012_out0;
wire v$_3013_out0;
wire v$_3014_out0;
wire v$_3015_out0;
wire v$_3051_out0;
wire v$_3052_out0;
wire v$_3053_out0;
wire v$_3054_out0;
wire v$_3055_out0;
wire v$_3056_out0;
wire v$_3057_out0;
wire v$_3058_out0;
wire v$_3059_out0;
wire v$_3060_out0;
wire v$_3061_out0;
wire v$_3062_out0;
wire v$_3063_out0;
wire v$_3064_out0;
wire v$_3065_out0;
wire v$_3066_out0;
wire v$_3067_out0;
wire v$_3068_out0;
wire v$_3069_out0;
wire v$_3070_out0;
wire v$_3071_out0;
wire v$_3072_out0;
wire v$_3073_out0;
wire v$_3074_out0;
wire v$_3075_out0;
wire v$_3076_out0;
wire v$_3077_out0;
wire v$_3078_out0;
wire v$_3079_out0;
wire v$_3080_out0;
wire v$_3085_out0;
wire v$_3086_out0;
wire v$_3087_out0;
wire v$_3088_out0;
wire v$_3089_out0;
wire v$_3090_out0;
wire v$_3091_out0;
wire v$_3092_out0;
wire v$_3093_out0;
wire v$_3094_out0;
wire v$_3095_out0;
wire v$_3096_out0;
wire v$_3097_out0;
wire v$_3098_out0;
wire v$_3099_out0;
wire v$_3100_out0;
wire v$_3101_out0;
wire v$_3102_out0;
wire v$_3103_out0;
wire v$_3104_out0;
wire v$_3105_out0;
wire v$_3106_out0;
wire v$_3107_out0;
wire v$_3108_out0;
wire v$_3109_out0;
wire v$_3110_out0;
wire v$_3111_out0;
wire v$_3112_out0;
wire v$_3113_out0;
wire v$_3114_out0;
wire v$_3119_out0;
wire v$_3120_out0;
wire v$_3121_out0;
wire v$_3122_out0;
wire v$_3123_out0;
wire v$_3124_out0;
wire v$_3139_out0;
wire v$_3140_out0;
wire v$_3141_out0;
wire v$_3142_out0;
wire v$_3143_out0;
wire v$_3144_out0;
wire v$_3145_out0;
wire v$_3146_out0;
wire v$_3147_out0;
wire v$_3148_out0;
wire v$_3149_out0;
wire v$_3150_out0;
wire v$_3151_out0;
wire v$_3152_out0;
wire v$_3153_out0;
wire v$_3154_out0;
wire v$_3155_out0;
wire v$_3156_out0;
wire v$_3157_out0;
wire v$_3158_out0;
wire v$_3159_out0;
wire v$_3160_out0;
wire v$_3161_out0;
wire v$_3162_out0;
wire v$_3163_out0;
wire v$_3164_out0;
wire v$_3165_out0;
wire v$_3166_out0;
wire v$_3167_out0;
wire v$_3168_out0;
wire v$_3180_out0;
wire v$_3181_out0;
wire v$_3199_out0;
wire v$_3200_out0;
wire v$_321_out0;
wire v$_322_out0;
wire v$_3237_out0;
wire v$_3238_out0;
wire v$_323_out0;
wire v$_3247_out0;
wire v$_3248_out0;
wire v$_3249_out0;
wire v$_324_out0;
wire v$_3250_out0;
wire v$_3266_out0;
wire v$_3267_out0;
wire v$_3270_out0;
wire v$_3271_out0;
wire v$_3282_out0;
wire v$_3283_out0;
wire v$_3284_out0;
wire v$_3285_out0;
wire v$_329_out0;
wire v$_330_out0;
wire v$_331_out0;
wire v$_332_out0;
wire v$_37_out0;
wire v$_3803_out0;
wire v$_3804_out0;
wire v$_3823_out0;
wire v$_3824_out0;
wire v$_3825_out0;
wire v$_3826_out0;
wire v$_3827_out0;
wire v$_3828_out0;
wire v$_3829_out0;
wire v$_3830_out0;
wire v$_3831_out0;
wire v$_3832_out0;
wire v$_3833_out0;
wire v$_3834_out0;
wire v$_3835_out0;
wire v$_3836_out0;
wire v$_3837_out0;
wire v$_3838_out0;
wire v$_3839_out0;
wire v$_3840_out0;
wire v$_3841_out0;
wire v$_3842_out0;
wire v$_3843_out0;
wire v$_3844_out0;
wire v$_3845_out0;
wire v$_3846_out0;
wire v$_3847_out0;
wire v$_3848_out0;
wire v$_3849_out0;
wire v$_3850_out0;
wire v$_3851_out0;
wire v$_3852_out0;
wire v$_3861_out0;
wire v$_3862_out0;
wire v$_3863_out0;
wire v$_3864_out0;
wire v$_3865_out0;
wire v$_3866_out0;
wire v$_3867_out0;
wire v$_3868_out0;
wire v$_3869_out0;
wire v$_3870_out0;
wire v$_3871_out0;
wire v$_3872_out0;
wire v$_3873_out0;
wire v$_3874_out0;
wire v$_3875_out0;
wire v$_3876_out0;
wire v$_3877_out0;
wire v$_3878_out0;
wire v$_3879_out0;
wire v$_3880_out0;
wire v$_3881_out0;
wire v$_3882_out0;
wire v$_3883_out0;
wire v$_3884_out0;
wire v$_3885_out0;
wire v$_3886_out0;
wire v$_3887_out0;
wire v$_3888_out0;
wire v$_3889_out0;
wire v$_3890_out0;
wire v$_38_out0;
wire v$_3907_out0;
wire v$_3908_out0;
wire v$_3910_out0;
wire v$_3911_out0;
wire v$_3912_out0;
wire v$_3913_out0;
wire v$_3914_out0;
wire v$_3915_out0;
wire v$_3916_out0;
wire v$_3917_out0;
wire v$_3918_out0;
wire v$_3919_out0;
wire v$_3920_out0;
wire v$_3921_out0;
wire v$_3922_out0;
wire v$_3923_out0;
wire v$_3924_out0;
wire v$_3925_out0;
wire v$_3926_out0;
wire v$_3927_out0;
wire v$_3928_out0;
wire v$_3929_out0;
wire v$_3930_out0;
wire v$_3931_out0;
wire v$_3932_out0;
wire v$_3933_out0;
wire v$_3934_out0;
wire v$_3935_out0;
wire v$_3936_out0;
wire v$_3937_out0;
wire v$_3938_out0;
wire v$_3939_out0;
wire v$_3961_out0;
wire v$_3962_out0;
wire v$_3963_out0;
wire v$_3964_out0;
wire v$_3965_out0;
wire v$_3966_out0;
wire v$_3967_out0;
wire v$_3968_out0;
wire v$_3969_out0;
wire v$_3970_out0;
wire v$_3971_out0;
wire v$_3972_out0;
wire v$_3973_out0;
wire v$_3974_out0;
wire v$_3975_out0;
wire v$_3976_out0;
wire v$_3977_out0;
wire v$_3978_out0;
wire v$_3979_out0;
wire v$_3980_out0;
wire v$_3981_out0;
wire v$_3982_out0;
wire v$_3983_out0;
wire v$_3984_out0;
wire v$_3985_out0;
wire v$_3986_out0;
wire v$_3987_out0;
wire v$_3988_out0;
wire v$_3989_out0;
wire v$_3990_out0;
wire v$_3_out0;
wire v$_413_out0;
wire v$_414_out0;
wire v$_437_out0;
wire v$_438_out0;
wire v$_4526_out1;
wire v$_4527_out1;
wire v$_4597_out0;
wire v$_4598_out0;
wire v$_4599_out0;
wire v$_4600_out0;
wire v$_4605_out0;
wire v$_4605_out1;
wire v$_4606_out0;
wire v$_4606_out1;
wire v$_4610_out0;
wire v$_4611_out0;
wire v$_468_out0;
wire v$_469_out0;
wire v$_470_out0;
wire v$_4711_out0;
wire v$_4712_out0;
wire v$_4713_out0;
wire v$_4714_out0;
wire v$_471_out0;
wire v$_472_out0;
wire v$_473_out0;
wire v$_474_out0;
wire v$_475_out0;
wire v$_476_out0;
wire v$_477_out0;
wire v$_478_out0;
wire v$_479_out0;
wire v$_480_out0;
wire v$_4812_out0;
wire v$_4813_out0;
wire v$_4814_out0;
wire v$_4815_out0;
wire v$_481_out0;
wire v$_482_out0;
wire v$_4831_out1;
wire v$_4832_out1;
wire v$_4833_out0;
wire v$_4834_out0;
wire v$_4837_out0;
wire v$_4838_out0;
wire v$_483_out0;
wire v$_484_out0;
wire v$_4856_out0;
wire v$_4857_out0;
wire v$_485_out0;
wire v$_486_out0;
wire v$_487_out0;
wire v$_488_out0;
wire v$_489_out0;
wire v$_490_out0;
wire v$_491_out0;
wire v$_492_out0;
wire v$_493_out0;
wire v$_494_out0;
wire v$_495_out0;
wire v$_496_out0;
wire v$_497_out0;
wire v$_503_out0;
wire v$_504_out0;
wire v$_505_out0;
wire v$_506_out0;
wire v$_507_out0;
wire v$_508_out0;
wire v$_509_out0;
wire v$_510_out0;
wire v$_511_out0;
wire v$_512_out0;
wire v$_513_out0;
wire v$_514_out0;
wire v$_515_out0;
wire v$_516_out0;
wire v$_517_out0;
wire v$_518_out0;
wire v$_519_out0;
wire v$_520_out0;
wire v$_521_out0;
wire v$_522_out0;
wire v$_523_out0;
wire v$_524_out0;
wire v$_525_out0;
wire v$_526_out0;
wire v$_527_out0;
wire v$_528_out0;
wire v$_529_out0;
wire v$_530_out0;
wire v$_531_out0;
wire v$_532_out0;
wire v$_568_out0;
wire v$_569_out0;
wire v$_570_out0;
wire v$_571_out0;
wire v$_572_out0;
wire v$_573_out0;
wire v$_574_out0;
wire v$_575_out0;
wire v$_576_out0;
wire v$_577_out0;
wire v$_578_out0;
wire v$_579_out0;
wire v$_580_out0;
wire v$_581_out0;
wire v$_582_out0;
wire v$_5832_out0;
wire v$_5832_out1;
wire v$_5833_out0;
wire v$_5833_out1;
wire v$_583_out0;
wire v$_584_out0;
wire v$_585_out0;
wire v$_5860_out0;
wire v$_5860_out1;
wire v$_586_out0;
wire v$_587_out0;
wire v$_588_out0;
wire v$_589_out0;
wire v$_590_out0;
wire v$_591_out0;
wire v$_592_out0;
wire v$_593_out0;
wire v$_594_out0;
wire v$_595_out0;
wire v$_596_out0;
wire v$_597_out0;
wire v$_60_out0;
wire v$_61_out0;
wire v$_6800_out0;
wire v$_6801_out0;
wire v$_6802_out0;
wire v$_6803_out0;
wire v$_6804_out0;
wire v$_6805_out0;
wire v$_6806_out0;
wire v$_6807_out0;
wire v$_6808_out0;
wire v$_6809_out0;
wire v$_6810_out0;
wire v$_6811_out0;
wire v$_6812_out0;
wire v$_6813_out0;
wire v$_6814_out0;
wire v$_6815_out0;
wire v$_6816_out0;
wire v$_6817_out0;
wire v$_6818_out0;
wire v$_6819_out0;
wire v$_6820_out0;
wire v$_6821_out0;
wire v$_6822_out0;
wire v$_6823_out0;
wire v$_6824_out0;
wire v$_6825_out0;
wire v$_6826_out0;
wire v$_6827_out0;
wire v$_6828_out0;
wire v$_6829_out0;
wire v$_6830_out0;
wire v$_6831_out0;
wire v$_6832_out0;
wire v$_6833_out0;
wire v$_6834_out0;
wire v$_6835_out0;
wire v$_6836_out0;
wire v$_6837_out0;
wire v$_6838_out0;
wire v$_6839_out0;
wire v$_6840_out0;
wire v$_6841_out0;
wire v$_6842_out0;
wire v$_6843_out0;
wire v$_6844_out0;
wire v$_6845_out0;
wire v$_6846_out0;
wire v$_6847_out0;
wire v$_6848_out0;
wire v$_6849_out0;
wire v$_6850_out0;
wire v$_6851_out0;
wire v$_6852_out0;
wire v$_6853_out0;
wire v$_6854_out0;
wire v$_6855_out0;
wire v$_6856_out0;
wire v$_6857_out0;
wire v$_6858_out0;
wire v$_6859_out0;
wire v$_6876_out0;
wire v$_6876_out1;
wire v$_6877_out0;
wire v$_6877_out1;
wire v$_7062_out1;
wire v$_7063_out1;
wire v$_7070_out0;
wire v$_7071_out0;
wire v$_7095_out0;
wire v$_7096_out0;
wire v$_7108_out0;
wire v$_7109_out0;
wire v$_7644_out0;
wire v$_7645_out0;
wire v$_7646_out0;
wire v$_7647_out0;
wire v$_7648_out0;
wire v$_7649_out0;
wire v$_7650_out0;
wire v$_7651_out0;
wire v$_7652_out0;
wire v$_7653_out0;
wire v$_7654_out0;
wire v$_7655_out0;
wire v$_7656_out0;
wire v$_7657_out0;
wire v$_7658_out0;
wire v$_7659_out0;
wire v$_7660_out0;
wire v$_7661_out0;
wire v$_7662_out0;
wire v$_7663_out0;
wire v$_7664_out0;
wire v$_7665_out0;
wire v$_7666_out0;
wire v$_7667_out0;
wire v$_7668_out0;
wire v$_7669_out0;
wire v$_7670_out0;
wire v$_7671_out0;
wire v$_7672_out0;
wire v$_7673_out0;
wire v$_77_out0;
wire v$_78_out0;
wire v$_79_out0;
wire v$_80_out0;
wire v$_8699_out0;
wire v$_8700_out0;
wire v$_8701_out0;
wire v$_8702_out0;
wire v$_8703_out0;
wire v$_8704_out0;
wire v$_8705_out0;
wire v$_8706_out0;
wire v$_8707_out0;
wire v$_8708_out0;
wire v$_8709_out0;
wire v$_8710_out0;
wire v$_8711_out0;
wire v$_8712_out0;
wire v$_8713_out0;
wire v$_8714_out0;
wire v$_8715_out0;
wire v$_8716_out0;
wire v$_8717_out0;
wire v$_8718_out0;
wire v$_8719_out0;
wire v$_8720_out0;
wire v$_8721_out0;
wire v$_8722_out0;
wire v$_8723_out0;
wire v$_8724_out0;
wire v$_8725_out0;
wire v$_8726_out0;
wire v$_8727_out0;
wire v$_8728_out0;
wire v$_8748_out0;
wire v$_8749_out0;
wire v$_8750_out0;
wire v$_8751_out0;
wire v$_8769_out0;
wire v$_8770_out0;
wire v$_8771_out0;
wire v$_8772_out0;
wire v$_8773_out0;
wire v$_8774_out0;
wire v$_8775_out0;
wire v$_8776_out0;
wire v$_8777_out0;
wire v$_8778_out0;
wire v$_8779_out0;
wire v$_8780_out0;
wire v$_8781_out0;
wire v$_8782_out0;
wire v$_8783_out0;
wire v$_8784_out0;
wire v$_8785_out0;
wire v$_8786_out0;
wire v$_8787_out0;
wire v$_8788_out0;
wire v$_8789_out0;
wire v$_8790_out0;
wire v$_8791_out0;
wire v$_8792_out0;
wire v$_8793_out0;
wire v$_8794_out0;
wire v$_8795_out0;
wire v$_8796_out0;
wire v$_8797_out0;
wire v$_8798_out0;
wire v$_8827_out0;
wire v$_8828_out0;
wire v$_8829_out0;
wire v$_8830_out0;
wire v$_8831_out0;
wire v$_8832_out0;
wire v$_8848_out0;
wire v$_8849_out0;
wire v$_8850_out0;
wire v$_8851_out0;
wire v$byte$comp$10_2318_out0;
wire v$byte$comp$11_2645_out0;
wire v$byte$comp$1_6872_out0;
wire v$byte$comp$1_6923_out0;
wire v$byte$ready_5842_out0;
wire v$byte$ready_5843_out0;
wire v$done$receiving_10604_out0;
wire v$exec1ls_3341_out0;
wire v$exec1ls_3342_out0;
wire v$transmit$INSTRUCTION_2674_out0;
wire v$wen$ram_4595_out0;
wire v$wen$ram_4596_out0;

always @(posedge clk) v$FF1_48_out0 <= v$BYTE$READY_2852_out0;
always @(posedge clk) v$FF1_49_out0 <= v$BYTE$READY_2853_out0;
always @(posedge clk) v$FF6_112_out0 <= v$ENABLE_2651_out0 ? v$MUX5_13348_out0 : v$FF6_112_out0;
always @(posedge clk) v$REG1_432_out0 <= v$G19_10327_out0 ? v$MUX4_2658_out0 : v$REG1_432_out0;
always @(posedge clk) v$REG1_433_out0 <= v$G19_10328_out0 ? v$MUX4_2659_out0 : v$REG1_433_out0;
v$ROM1_462 I462 (v$ROM1_462_out0, v$REG1_7134_out0, clk);
always @(posedge clk) v$FF4_463_out0 <= v$ENABLE_2651_out0 ? v$MUX3_7140_out0 : v$FF4_463_out0;
v$RAM0_1680 I1680 (v$RAM0_1680_out0, v$ADRESS$ins0_11169_out0, v$DATA$RAM$IN0_284_out0, v$DONE$RECEIVING_5857_out0, clk);
v$data$ram_1818 I1818 (v$data$ram_1818_out0, v$ADRESS_8683_out0, v$DATA_2469_out0, v$WEN_2154_out0, clk);
always @(posedge clk) v$FF1_1955_out0 <= v$ENABLE_2651_out0 ? v$SEL1_13445_out0 : v$FF1_1955_out0;
always @(posedge clk) v$IHOLD$REGISTER_2013_out0 <= v$NORMAL_181_out0 ? v$RAM$OUT_1751_out0 : v$IHOLD$REGISTER_2013_out0;
always @(posedge clk) v$IHOLD$REGISTER_2014_out0 <= v$NORMAL_182_out0 ? v$RAM$OUT_1752_out0 : v$IHOLD$REGISTER_2014_out0;
always @(posedge clk) v$FF3_2016_out0 <= v$EN_7093_out0 ? v$_4605_out0 : v$FF3_2016_out0;
always @(posedge clk) v$FF3_2017_out0 <= v$EN_7094_out0 ? v$_4606_out0 : v$FF3_2017_out0;
always @(posedge clk) v$FF4_2106_out0 <= v$EN_7093_out0 ? v$_4605_out1 : v$FF4_2106_out0;
always @(posedge clk) v$FF4_2107_out0 <= v$EN_7094_out0 ? v$_4606_out1 : v$FF4_2107_out0;
always @(posedge clk) v$REG1_2314_out0 <= v$D1_8842_out1 ? v$DIN3_10310_out0 : v$REG1_2314_out0;
always @(posedge clk) v$REG1_2315_out0 <= v$D1_8843_out1 ? v$DIN3_10311_out0 : v$REG1_2315_out0;
always @(posedge clk) v$FF7_2670_out0 <= v$G24_10560_out0;
always @(posedge clk) v$FF7_2671_out0 <= v$G24_10561_out0;
always @(posedge clk) v$FF7_2672_out0 <= v$G24_10562_out0;
always @(posedge clk) v$FF7_2673_out0 <= v$G24_10563_out0;
always @(posedge clk) v$REG1_2677_out0 <= v$ENABLE_1757_out0 ? v$_3040_out0 : v$REG1_2677_out0;
always @(posedge clk) v$FF2_2833_out0 <= v$ENABLE_2651_out0 ? v$MUX1_2625_out0 : v$FF2_2833_out0;
always @(posedge clk) v$FF1_4717_out0 <= v$EN_2919_out0 ? v$G1_2700_out0 : v$FF1_4717_out0;
always @(posedge clk) v$FF1_4718_out0 <= v$EN_2920_out0 ? v$G1_2701_out0 : v$FF1_4718_out0;
always @(posedge clk) v$FF1_4719_out0 <= v$EN_2921_out0 ? v$G1_2702_out0 : v$FF1_4719_out0;
always @(posedge clk) v$FF1_4720_out0 <= v$EN_2922_out0 ? v$G1_2703_out0 : v$FF1_4720_out0;
always @(posedge clk) v$FF1_4721_out0 <= v$EN_2923_out0 ? v$G1_2704_out0 : v$FF1_4721_out0;
always @(posedge clk) v$FF1_4722_out0 <= v$EN_2924_out0 ? v$G1_2705_out0 : v$FF1_4722_out0;
always @(posedge clk) v$FF1_4723_out0 <= v$EN_2925_out0 ? v$G1_2706_out0 : v$FF1_4723_out0;
always @(posedge clk) v$FF1_4724_out0 <= v$EN_2926_out0 ? v$G1_2707_out0 : v$FF1_4724_out0;
always @(posedge clk) v$FF1_4725_out0 <= v$EN_2927_out0 ? v$G1_2708_out0 : v$FF1_4725_out0;
always @(posedge clk) v$FF1_4726_out0 <= v$EN_2928_out0 ? v$G1_2709_out0 : v$FF1_4726_out0;
always @(posedge clk) v$FF1_4727_out0 <= v$EN_2929_out0 ? v$G1_2710_out0 : v$FF1_4727_out0;
always @(posedge clk) v$FF1_4728_out0 <= v$EN_2930_out0 ? v$G1_2711_out0 : v$FF1_4728_out0;
always @(posedge clk) v$FF1_4729_out0 <= v$EN_2931_out0 ? v$G1_2712_out0 : v$FF1_4729_out0;
always @(posedge clk) v$FF1_4730_out0 <= v$EN_2932_out0 ? v$G1_2713_out0 : v$FF1_4730_out0;
always @(posedge clk) v$FF1_4731_out0 <= v$EN_2933_out0 ? v$G1_2714_out0 : v$FF1_4731_out0;
always @(posedge clk) v$FF1_4732_out0 <= v$EN_2934_out0 ? v$G1_2715_out0 : v$FF1_4732_out0;
always @(posedge clk) v$REG3_4747_out0 <= v$D1_8842_out3 ? v$DIN3_10310_out0 : v$REG3_4747_out0;
always @(posedge clk) v$REG3_4748_out0 <= v$D1_8843_out3 ? v$DIN3_10311_out0 : v$REG3_4748_out0;
always @(posedge clk) v$FF7_4781_out0 <= v$ENABLE_2651_out0 ? v$MUX6_10976_out0 : v$FF7_4781_out0;
always @(posedge clk) v$FF1_4841_out0 <= v$G20_11040_out0;
always @(posedge clk) v$REG1_7031_out0 <= v$G8_7103_out0 ? v$MUX1_11061_out0 : v$REG1_7031_out0;
always @(posedge clk) v$FF5_7100_out0 <= v$ENABLE_2651_out0 ? v$MUX4_3219_out0 : v$FF5_7100_out0;
always @(posedge clk) v$REG1_7134_out0 <= v$EQ3_5861_out0 ? v$A1_11043_out0 : v$REG1_7134_out0;
always @(posedge clk) v$FF9_8805_out0 <= v$ENABLE_2651_out0 ? v$MUX8_2697_out0 : v$FF9_8805_out0;
always @(posedge clk) v$FF1_10325_out0 <= v$G3_2941_out0 ? v$G2_10799_out0 : v$FF1_10325_out0;
always @(posedge clk) v$FF1_10326_out0 <= v$G3_2942_out0 ? v$G2_10800_out0 : v$FF1_10326_out0;
always @(posedge clk) v$REG1_10368_out0 <= v$_533_out0;
always @(posedge clk) v$REG1_10546_out0 <= v$G8_16_out0 ? v$OUT_3037_out0 : v$REG1_10546_out0;
always @(posedge clk) v$FF8_10849_out0 <= v$G21_3808_out0;
always @(posedge clk) v$FF8_10850_out0 <= v$G21_3809_out0;
always @(posedge clk) v$FF8_10851_out0 <= v$G21_3810_out0;
always @(posedge clk) v$FF8_10852_out0 <= v$G21_3811_out0;
always @(posedge clk) v$REG0_10912_out0 <= v$D1_8842_out0 ? v$DIN3_10310_out0 : v$REG0_10912_out0;
always @(posedge clk) v$REG0_10913_out0 <= v$D1_8843_out0 ? v$DIN3_10311_out0 : v$REG0_10913_out0;
always @(posedge clk) v$FF3_11046_out0 <= v$ENABLE_2651_out0 ? v$MUX2_4448_out0 : v$FF3_11046_out0;
always @(posedge clk) v$FF2_11062_out0 <= v$FF1_13511_out0;
always @(posedge clk) v$REG1_11130_out0 <= v$G2_6884_out0 ? v$COUT_3895_out0 : v$REG1_11130_out0;
always @(posedge clk) v$REG1_11131_out0 <= v$G2_6885_out0 ? v$COUT_3896_out0 : v$REG1_11131_out0;
always @(posedge clk) v$FF8_11222_out0 <= v$ENABLE_2651_out0 ? v$MUX7_10448_out0 : v$FF8_11222_out0;
always @(posedge clk) v$REG2_12251_out0 <= v$D1_8842_out2 ? v$DIN3_10310_out0 : v$REG2_12251_out0;
always @(posedge clk) v$REG2_12252_out0 <= v$D1_8843_out2 ? v$DIN3_10311_out0 : v$REG2_12252_out0;
always @(posedge clk) v$REG1_13338_out0 <= v$COUT_10922_out0;
always @(posedge clk) v$REG1_13339_out0 <= v$COUT_10937_out0;
v$RAM1_13398 I13398 (v$RAM1_13398_out0, v$ADRESS$ins1_10617_out0, v$DATA$RAM$IN1_4779_out0, v$C3_2764_out0, clk);
always @(posedge clk) v$FF1_13511_out0 <= v$ROM1_462_out0;
assign v$C11_13766_out0 = 6'h0;
assign v$C11_13765_out0 = 6'h0;
assign v$C1_13447_out0 = 8'h0;
assign v$C1_13446_out0 = 8'h0;
assign v$C1_13278_out0 = 8'h0;
assign v$C1_13277_out0 = 8'h0;
assign v$C5_13267_out0 = 1'h1;
assign v$C1_11293_out0 = 2'h0;
assign v$C1_11292_out0 = 2'h0;
assign v$C10_11249_out0 = 5'h1f;
assign v$C10_11248_out0 = 5'h1f;
assign v$C2_11233_out0 = 3'h0;
assign v$C9_11160_out0 = 6'h3f;
assign v$C9_11159_out0 = 6'h3f;
assign v$C5_11031_out0 = 1'h0;
assign v$C3_10853_out0 = 3'h0;
assign v$C14_10796_out0 = 5'h1;
assign v$C14_10795_out0 = 5'h1;
assign v$C1_10790_out0 = 1'h0;
assign v$C1_10789_out0 = 1'h0;
assign v$C2_10762_out0 = 12'h7ff;
assign v$C2_10761_out0 = 12'h7ff;
assign v$C4_10619_out0 = 1'h1;
assign v$C5_10356_out0 = 2'h0;
assign v$C6_10318_out0 = 1'h1;
assign v$C6_10317_out0 = 1'h1;
assign v$C1_10316_out0 = 5'h0;
assign v$C1_10315_out0 = 5'h0;
assign v$C1_10314_out0 = 5'h0;
assign v$C1_10313_out0 = 5'h0;
assign v$C1_10306_out0 = 4'h0;
assign v$C1_10305_out0 = 4'h0;
assign v$C1_10267_out0 = 8'h0;
assign v$C1_10266_out0 = 8'h0;
assign v$C1_10259_out0 = 1'h0;
assign v$C1_8816_out0 = 1'h0;
assign v$C1_8815_out0 = 1'h0;
assign v$2_7072_out0 = 1'h1;
assign v$C1_6920_out0 = 4'h0;
assign v$C1_6919_out0 = 4'h0;
assign v$C1_6794_out0 = 2'h0;
assign v$C1_6793_out0 = 2'h0;
assign v$C3_4742_out0 = 1'h0;
assign v$C3_4741_out0 = 1'h0;
assign v$C11_4540_out0 = 16'hffff;
assign v$C11_4539_out0 = 16'hffff;
assign v$C7_3222_out0 = 1'h1;
assign v$C1_3211_out0 = 12'h0;
assign v$C1_3210_out0 = 12'h0;
assign v$C1_3206_out0 = 2'h0;
assign v$C1_3205_out0 = 2'h0;
assign v$C9_3030_out0 = 1'h0;
assign v$C9_3029_out0 = 1'h0;
assign v$C3_2764_out0 = 1'h0;
assign v$C8_2759_out0 = 5'h0;
assign v$C8_2758_out0 = 5'h0;
assign v$C1_2716_out0 = 3'h0;
assign v$C5_2689_out0 = 16'hffff;
assign v$C5_2688_out0 = 16'hffff;
assign v$C4_2594_out0 = 5'h0;
assign v$C4_2593_out0 = 5'h0;
assign v$C1_2427_out0 = 12'h7f4;
assign v$C1_2426_out0 = 12'h7f4;
assign v$C2_2413_out0 = 12'h0;
assign v$C7_2272_out0 = 1'h0;
assign v$C7_2271_out0 = 1'h0;
assign v$C13_2186_out0 = 16'h0;
assign v$C13_2185_out0 = 16'h0;
assign v$C12_2114_out0 = 6'hf;
assign v$C12_2113_out0 = 6'hf;
assign v$C1_2006_out0 = 4'h4;
assign v$C1_2005_out0 = 4'h4;
assign v$C7_1866_out0 = 16'h0;
assign v$C7_1865_out0 = 16'h0;
assign v$C10_1820_out0 = 1'h1;
assign v$C10_1819_out0 = 1'h1;
assign v$C_1808_out0 = 11'h0;
assign v$C_1807_out0 = 11'h0;
assign v$C6_1732_out0 = 1'h1;
assign v$C15_1731_out0 = 16'hffff;
assign v$C15_1730_out0 = 16'hffff;
assign v$C14_1675_out0 = 1'h1;
assign v$C14_1674_out0 = 1'h1;
assign v$C4_1201_out0 = 3'h0;
assign v$C12_1152_out0 = 1'h1;
assign v$C12_1151_out0 = 1'h1;
assign v$C1_607_out0 = 11'h0;
assign v$C1_606_out0 = 11'h0;
assign v$C1_605_out0 = 1'h0;
assign v$C1_604_out0 = 1'h0;
assign v$C1_436_out0 = 1'h1;
assign v$C13_406_out0 = 6'h31;
assign v$C13_405_out0 = 6'h31;
assign v$C4_90_out0 = 1'h0;
assign v$ROR_67_out0 = 2'h3;
assign v$ROR_66_out0 = 2'h3;
assign v$Q_291_out0 = v$FF1_4717_out0;
assign v$Q_292_out0 = v$FF1_4718_out0;
assign v$Q_293_out0 = v$FF1_4719_out0;
assign v$Q_294_out0 = v$FF1_4720_out0;
assign v$Q_295_out0 = v$FF1_4721_out0;
assign v$Q_296_out0 = v$FF1_4722_out0;
assign v$Q_297_out0 = v$FF1_4723_out0;
assign v$Q_298_out0 = v$FF1_4724_out0;
assign v$Q_299_out0 = v$FF1_4725_out0;
assign v$Q_300_out0 = v$FF1_4726_out0;
assign v$Q_301_out0 = v$FF1_4727_out0;
assign v$Q_302_out0 = v$FF1_4728_out0;
assign v$Q_303_out0 = v$FF1_4729_out0;
assign v$Q_304_out0 = v$FF1_4730_out0;
assign v$Q_305_out0 = v$FF1_4731_out0;
assign v$Q_306_out0 = v$FF1_4732_out0;
assign v$DATA$OUT_1135_out0 = v$data$ram_1818_out0;
assign v$EQ4_1142_out0 = v$REG1_7134_out0 == 12'h0;
assign v$_1673_out0 = { v$FF1_4841_out0,v$C2_11233_out0 };
assign v$R0_1688_out0 = v$REG0_10912_out0;
assign v$R0_1689_out0 = v$REG0_10913_out0;
assign v$Q6_1889_out0 = v$FF7_2670_out0;
assign v$Q6_1890_out0 = v$FF7_2671_out0;
assign v$Q6_1891_out0 = v$FF7_2672_out0;
assign v$Q6_1892_out0 = v$FF7_2673_out0;
assign v$DIV$INST_2324_out0 = v$DIV$INST1_7011_out0;
assign v$DIV$INST_2325_out0 = v$DIV$INST0_6905_out0;
assign v$RAM$OUT1_2385_out0 = v$RAM1_13398_out0;
assign v$IR_2826_out0 = v$IHOLD$REGISTER_2013_out0;
assign v$IR_2827_out0 = v$IHOLD$REGISTER_2014_out0;
assign v$_2887_out0 = { v$FF3_2016_out0,v$FF4_2106_out0 };
assign v$_2888_out0 = { v$FF3_2017_out0,v$FF4_2107_out0 };
assign v$_2959_out0 = v$REG1_2677_out0[0:0];
assign v$_2959_out1 = v$REG1_2677_out0[7:7];
assign v$OUT_3037_out0 = v$REG1_2677_out0;
assign v$R2_3043_out0 = v$REG2_12251_out0;
assign v$R2_3044_out0 = v$REG2_12252_out0;
assign v$C_3197_out0 = v$REG1_11130_out0;
assign v$C_3198_out0 = v$REG1_11131_out0;
assign v$C_3207_out0 = v$REG1_11130_out0;
assign v$C_3208_out0 = v$REG1_11131_out0;
assign v$EQ1_3344_out0 = v$REG1_7031_out0 == 2'h2;
assign v$Q1_3993_out0 = v$FF1_4841_out0;
assign v$EN_4485_out0 = v$C5_13267_out0;
assign v$R3_4652_out0 = v$REG3_4747_out0;
assign v$R3_4653_out0 = v$REG3_4748_out0;
assign v$byte$ready_5842_out0 = v$C5_11031_out0;
assign v$_5860_out0 = v$REG1_10368_out0[0:0];
assign v$_5860_out1 = v$REG1_10368_out0[1:1];
assign v$Q7_6888_out0 = v$FF8_10849_out0;
assign v$Q7_6889_out0 = v$FF8_10850_out0;
assign v$Q7_6890_out0 = v$FF8_10851_out0;
assign v$Q7_6891_out0 = v$FF8_10852_out0;
assign v$NEG1_6921_out0 = v$C9_11159_out0;
assign v$NEG1_6922_out0 = v$C9_11160_out0;
assign v$_7116_out0 = v$IHOLD$REGISTER_2013_out0[11:0];
assign v$_7116_out1 = v$IHOLD$REGISTER_2013_out0[15:4];
assign v$_7117_out0 = v$IHOLD$REGISTER_2014_out0[11:0];
assign v$_7117_out1 = v$IHOLD$REGISTER_2014_out0[15:4];
assign v$RECEIVERSTREAM_7635_out0 = v$REG1_10546_out0;
assign v$RX$BYTEREADY_8756_out0 = v$FF1_4841_out0;
assign v$R1_8761_out0 = v$REG1_2314_out0;
assign v$R1_8762_out0 = v$REG1_2315_out0;
assign v$RAM$OUT0_8764_out0 = v$RAM0_1680_out0;
assign v$0B00001_10554_out0 = v$C14_10795_out0;
assign v$0B00001_10555_out0 = v$C14_10796_out0;
assign v$Q_10618_out0 = v$REG1_10368_out0;
assign v$0_10706_out0 = v$C7_2271_out0;
assign v$0_10707_out0 = v$C7_2272_out0;
assign v$G2_10799_out0 = ! v$FF1_10325_out0;
assign v$G2_10800_out0 = ! v$FF1_10326_out0;
assign {v$A1_11043_out1,v$A1_11043_out0 } = v$C2_2413_out0 + v$REG1_7134_out0 + v$C1_436_out0;
assign v$FLOAT$INST16_13443_out0 = v$FF1_10325_out0;
assign v$FLOAT$INST16_13444_out0 = v$FF1_10326_out0;
assign v$Q_13510_out0 = v$REG1_7031_out0;
assign v$STALL$DUAL$CORE_13618_out0 = v$C4_90_out0;
assign v$SEL2_280_out0 = v$_7116_out0[9:9];
assign v$SEL2_281_out0 = v$_7117_out0[9:9];
assign v$MEM$RAM_434_out0 = v$DATA$OUT_1135_out0;
assign v$MEM$RAM_435_out0 = v$DATA$OUT_1135_out0;
assign v$RECEIVER$STREAM_564_out0 = v$RECEIVERSTREAM_7635_out0;
assign v$Q_1153_out0 = v$_2887_out0;
assign v$Q_1154_out0 = v$_2888_out0;
assign v$G5_1198_out0 = ! v$EN_4485_out0;
assign v$Q2_1676_out0 = v$Q_291_out0;
assign v$Q2_1677_out0 = v$Q_295_out0;
assign v$Q2_1678_out0 = v$Q_299_out0;
assign v$Q2_1679_out0 = v$Q_303_out0;
assign v$G10_1943_out0 = !(v$Q_292_out0 || v$Q_291_out0);
assign v$G10_1944_out0 = !(v$Q_296_out0 || v$Q_295_out0);
assign v$G10_1945_out0 = !(v$Q_300_out0 || v$Q_299_out0);
assign v$G10_1946_out0 = !(v$Q_304_out0 || v$Q_303_out0);
assign v$G4_1960_out0 = v$Q_294_out0 && v$Q_292_out0;
assign v$G4_1961_out0 = v$Q_298_out0 && v$Q_296_out0;
assign v$G4_1962_out0 = v$Q_302_out0 && v$Q_300_out0;
assign v$G4_1963_out0 = v$Q_306_out0 && v$Q_304_out0;
assign v$G28_2098_out0 = v$Q7_6888_out0 && v$Q6_1889_out0;
assign v$G28_2099_out0 = v$Q7_6889_out0 && v$Q6_1890_out0;
assign v$G28_2100_out0 = v$Q7_6890_out0 && v$Q6_1891_out0;
assign v$G28_2101_out0 = v$Q7_6891_out0 && v$Q6_1892_out0;
assign v$RAM$OUT_2104_out0 = v$RAM$OUT1_2385_out0;
assign v$RAM$OUT_2105_out0 = v$RAM$OUT0_8764_out0;
assign v$Q1_2112_out0 = v$_5860_out1;
assign v$EQ10_2320_out0 = v$_7116_out1 == 4'h3;
assign v$EQ10_2321_out0 = v$_7117_out1 == 4'h3;
assign v$RX$BYTE$READY_2436_out0 = v$RX$BYTEREADY_8756_out0;
assign v$_2536_out0 = { v$EQ1_3344_out0,v$C1_2716_out0 };
assign v$COUT_2725_out0 = v$A1_11043_out1;
assign v$R3TEST_2872_out0 = v$R3_4652_out0;
assign v$R3TEST_2873_out0 = v$R3_4653_out0;
assign v$FLOAT$INST_2955_out0 = v$FLOAT$INST16_13443_out0;
assign v$FLOAT$INST_2956_out0 = v$FLOAT$INST16_13444_out0;
assign v$G2_2975_out0 = ((v$Q_294_out0 && !v$Q_292_out0) || (!v$Q_294_out0) && v$Q_292_out0);
assign v$G2_2976_out0 = ((v$Q_298_out0 && !v$Q_296_out0) || (!v$Q_298_out0) && v$Q_296_out0);
assign v$G2_2977_out0 = ((v$Q_302_out0 && !v$Q_300_out0) || (!v$Q_302_out0) && v$Q_300_out0);
assign v$G2_2978_out0 = ((v$Q_306_out0 && !v$Q_304_out0) || (!v$Q_306_out0) && v$Q_304_out0);
assign v$_2983_out0 = v$Q_13510_out0[0:0];
assign v$_2983_out1 = v$Q_13510_out0[1:1];
assign v$R0TEST_3184_out0 = v$R0_1688_out0;
assign v$R0TEST_3185_out0 = v$R0_1689_out0;
assign v$G2_4468_out0 = ! v$STALL$DUAL$CORE_13618_out0;
assign v$NOTUSED_4609_out0 = v$_2959_out0;
assign v$EQ_4835_out0 = v$_7116_out1 == 4'h0;
assign v$EQ_4836_out0 = v$_7117_out1 == 4'h0;
assign v$G23_4852_out0 = ! v$Q7_6888_out0;
assign v$G23_4853_out0 = ! v$Q7_6889_out0;
assign v$G23_4854_out0 = ! v$Q7_6890_out0;
assign v$G23_4855_out0 = ! v$Q7_6891_out0;
assign v$RX$OVERFLOW_5848_out0 = v$EQ1_3344_out0;
assign v$EQ3_5861_out0 = v$Q_10618_out0 == 2'h3;
assign v$IR_7112_out0 = v$IR_2826_out0;
assign v$IR_7113_out0 = v$IR_2827_out0;
assign v$_7183_out0 = { v$Q7_6888_out0,v$Q6_1889_out0 };
assign v$_7184_out0 = { v$Q7_6889_out0,v$Q6_1890_out0 };
assign v$_7185_out0 = { v$Q7_6890_out0,v$Q6_1891_out0 };
assign v$_7186_out0 = { v$Q7_6891_out0,v$Q6_1892_out0 };
assign v$C_8648_out0 = v$C_3207_out0;
assign v$C_8649_out0 = v$C_3208_out0;
assign v$G1_8693_out0 = ! v$Q_294_out0;
assign v$G1_8694_out0 = ! v$Q_298_out0;
assign v$G1_8695_out0 = ! v$Q_302_out0;
assign v$G1_8696_out0 = ! v$Q_306_out0;
assign v$Q3_8737_out0 = v$Q_293_out0;
assign v$Q3_8738_out0 = v$Q_297_out0;
assign v$Q3_8739_out0 = v$Q_301_out0;
assign v$Q3_8740_out0 = v$Q_305_out0;
assign v$Q1_8859_out0 = v$Q_292_out0;
assign v$Q1_8860_out0 = v$Q_296_out0;
assign v$Q1_8861_out0 = v$Q_300_out0;
assign v$Q1_8862_out0 = v$Q_304_out0;
assign v$G9_10291_out0 = v$Q_294_out0 && v$Q_293_out0;
assign v$G9_10292_out0 = v$Q_298_out0 && v$Q_297_out0;
assign v$G9_10293_out0 = v$Q_302_out0 && v$Q_301_out0;
assign v$G9_10294_out0 = v$Q_306_out0 && v$Q_305_out0;
assign v$R1TEST_10485_out0 = v$R1_8761_out0;
assign v$R1TEST_10486_out0 = v$R1_8762_out0;
assign v$G24_10560_out0 = ((v$Q7_6888_out0 && !v$Q6_1889_out0) || (!v$Q7_6888_out0) && v$Q6_1889_out0);
assign v$G24_10561_out0 = ((v$Q7_6889_out0 && !v$Q6_1890_out0) || (!v$Q7_6889_out0) && v$Q6_1890_out0);
assign v$G24_10562_out0 = ((v$Q7_6890_out0 && !v$Q6_1891_out0) || (!v$Q7_6890_out0) && v$Q6_1891_out0);
assign v$G24_10563_out0 = ((v$Q7_6891_out0 && !v$Q6_1892_out0) || (!v$Q7_6891_out0) && v$Q6_1892_out0);
assign v$R2TEST_10708_out0 = v$R2_3043_out0;
assign v$R2TEST_10709_out0 = v$R2_3044_out0;
assign v$BYTE$READY_11172_out0 = v$byte$ready_5842_out0;
assign v$Q0_11198_out0 = v$Q_294_out0;
assign v$Q0_11199_out0 = v$Q_298_out0;
assign v$Q0_11200_out0 = v$Q_302_out0;
assign v$Q0_11201_out0 = v$Q_306_out0;
assign v$DIV$INSTRUCTION_11296_out0 = v$DIV$INST_2324_out0;
assign v$DIV$INSTRUCTION_11297_out0 = v$DIV$INST_2325_out0;
assign v$Q0_13351_out0 = v$_5860_out0;
assign v$NOUSED_13492_out0 = v$_7116_out0;
assign v$NOUSED_13493_out0 = v$_7117_out0;
assign v$EQ2_8_out0 = v$Q_1153_out0 == 2'h2;
assign v$EQ2_9_out0 = v$Q_1154_out0 == 2'h2;
assign v$R3TEST_117_out0 = v$R3TEST_2872_out0;
assign v$R3TEST_118_out0 = v$R3TEST_2873_out0;
assign v$LS_204_out0 = v$EQ_4835_out0;
assign v$LS_205_out0 = v$EQ_4836_out0;
assign v$4BITCOUNTER_317_out0 = v$_7183_out0;
assign v$4BITCOUNTER_318_out0 = v$_7184_out0;
assign v$4BITCOUNTER_319_out0 = v$_7185_out0;
assign v$4BITCOUNTER_320_out0 = v$_7186_out0;
assign v$EQ4_611_out0 = v$Q_1153_out0 == 2'h0;
assign v$EQ4_612_out0 = v$Q_1154_out0 == 2'h0;
assign v$G6_1159_out0 = v$G4_1960_out0 && v$Q_291_out0;
assign v$G6_1160_out0 = v$G4_1961_out0 && v$Q_295_out0;
assign v$G6_1161_out0 = v$G4_1962_out0 && v$Q_299_out0;
assign v$G6_1162_out0 = v$G4_1963_out0 && v$Q_303_out0;
assign v$IR_1871_out0 = v$IR_7112_out0;
assign v$IR_1872_out0 = v$IR_7113_out0;
assign v$G12_2270_out0 = ! v$Q1_2112_out0;
assign v$EQ1_2540_out0 = v$Q_1153_out0 == 2'h1;
assign v$EQ1_2541_out0 = v$Q_1154_out0 == 2'h1;
assign v$STALL$DUAL$CORE_3128_out0 = v$G2_4468_out0;
assign v$G3_3343_out0 = v$G5_1198_out0 && v$Q1_2112_out0;
assign v$G38_3903_out0 = v$Q2_1676_out0 || v$Q3_8737_out0;
assign v$G38_3904_out0 = v$Q2_1677_out0 || v$Q3_8738_out0;
assign v$G38_3905_out0 = v$Q2_1678_out0 || v$Q3_8739_out0;
assign v$G38_3906_out0 = v$Q2_1679_out0 || v$Q3_8740_out0;
assign v$RX$OVERFLOW_4469_out0 = v$RX$OVERFLOW_5848_out0;
assign v$Q0_4470_out0 = v$Q0_11198_out0;
assign v$Q0_4471_out0 = v$Q0_11199_out0;
assign v$Q0_4472_out0 = v$Q0_11200_out0;
assign v$Q0_4473_out0 = v$Q0_11201_out0;
assign v$G6_4818_out0 = ! v$_2983_out0;
assign v$C_4848_out0 = v$C_8648_out0;
assign v$C_4849_out0 = v$C_8649_out0;
assign v$_5832_out0 = v$Q_1153_out0[0:0];
assign v$_5832_out1 = v$Q_1153_out0[1:1];
assign v$_5833_out0 = v$Q_1154_out0[0:0];
assign v$_5833_out1 = v$Q_1154_out0[1:1];
assign v$Q2_6880_out0 = v$Q2_1676_out0;
assign v$Q2_6881_out0 = v$Q2_1677_out0;
assign v$Q2_6882_out0 = v$Q2_1678_out0;
assign v$Q2_6883_out0 = v$Q2_1679_out0;
assign v$G3_6894_out0 = ((v$G4_1960_out0 && !v$Q_291_out0) || (!v$G4_1960_out0) && v$Q_291_out0);
assign v$G3_6895_out0 = ((v$G4_1961_out0 && !v$Q_295_out0) || (!v$G4_1961_out0) && v$Q_295_out0);
assign v$G3_6896_out0 = ((v$G4_1962_out0 && !v$Q_299_out0) || (!v$G4_1962_out0) && v$Q_299_out0);
assign v$G3_6897_out0 = ((v$G4_1963_out0 && !v$Q_303_out0) || (!v$G4_1963_out0) && v$Q_303_out0);
assign v$G37_6900_out0 = v$Q1_8859_out0 || v$Q0_11198_out0;
assign v$G37_6901_out0 = v$Q1_8860_out0 || v$Q0_11199_out0;
assign v$G37_6902_out0 = v$Q1_8861_out0 || v$Q0_11200_out0;
assign v$G37_6903_out0 = v$Q1_8862_out0 || v$Q0_11201_out0;
assign v$Q1_6906_out0 = v$Q1_8859_out0;
assign v$Q1_6907_out0 = v$Q1_8860_out0;
assign v$Q1_6908_out0 = v$Q1_8861_out0;
assign v$Q1_6909_out0 = v$Q1_8862_out0;
assign v$G4_6914_out0 = ! v$Q0_13351_out0;
assign v$R0TEST_7005_out0 = v$R0TEST_3184_out0;
assign v$R0TEST_7006_out0 = v$R0TEST_3185_out0;
assign v$BYTE$READY_7021_out0 = v$BYTE$READY_11172_out0;
assign v$D_7680_out0 = v$G2_2975_out0;
assign v$D_7682_out0 = v$G1_8693_out0;
assign v$D_7684_out0 = v$G2_2976_out0;
assign v$D_7686_out0 = v$G1_8694_out0;
assign v$D_7688_out0 = v$G2_2977_out0;
assign v$D_7690_out0 = v$G1_8695_out0;
assign v$D_7692_out0 = v$G2_2978_out0;
assign v$D_7694_out0 = v$G1_8696_out0;
assign v$G11_8652_out0 = v$EN_4485_out0 && v$Q0_13351_out0;
assign v$G2_10278_out0 = ! v$EQ3_5861_out0;
assign v$RAM$OUT_10335_out0 = v$RAM$OUT_2104_out0;
assign v$RAM$OUT_10336_out0 = v$RAM$OUT_2105_out0;
assign v$_10376_out0 = { v$_1673_out0,v$_2536_out0 };
assign v$FLOATING$INSTRUCTION_10391_out0 = v$FLOAT$INST_2955_out0;
assign v$FLOATING$INSTRUCTION_10392_out0 = v$FLOAT$INST_2956_out0;
assign v$EN_10451_out0 = v$G28_2098_out0;
assign v$EN_10452_out0 = v$G28_2099_out0;
assign v$EN_10453_out0 = v$G28_2100_out0;
assign v$EN_10454_out0 = v$G28_2101_out0;
assign v$G1_10476_out0 = ! v$_2983_out1;
assign v$R1TEST_10498_out0 = v$R1TEST_10485_out0;
assign v$R1TEST_10499_out0 = v$R1TEST_10486_out0;
assign v$Q3_10518_out0 = v$Q3_8737_out0;
assign v$Q3_10519_out0 = v$Q3_8738_out0;
assign v$Q3_10520_out0 = v$Q3_8739_out0;
assign v$Q3_10521_out0 = v$Q3_8740_out0;
assign v$G8_10609_out0 = !(v$G9_10291_out0 && v$G10_1943_out0);
assign v$G8_10610_out0 = !(v$G9_10292_out0 && v$G10_1944_out0);
assign v$G8_10611_out0 = !(v$G9_10293_out0 && v$G10_1945_out0);
assign v$G8_10612_out0 = !(v$G9_10294_out0 && v$G10_1946_out0);
assign v$G8_10769_out0 = ! v$SEL2_280_out0;
assign v$G8_10770_out0 = ! v$SEL2_281_out0;
assign v$G1_10810_out0 = ((v$EN_4485_out0 && !v$Q0_13351_out0) || (!v$EN_4485_out0) && v$Q0_13351_out0);
assign v$G22_10983_out0 = v$G23_4852_out0 && v$Q6_1889_out0;
assign v$G22_10984_out0 = v$G23_4853_out0 && v$Q6_1890_out0;
assign v$G22_10985_out0 = v$G23_4854_out0 && v$Q6_1891_out0;
assign v$G22_10986_out0 = v$G23_4855_out0 && v$Q6_1892_out0;
assign v$R2TEST_10987_out0 = v$R2TEST_10708_out0;
assign v$R2TEST_10988_out0 = v$R2TEST_10709_out0;
assign v$RAM$OUT_11214_out0 = v$MEM$RAM_434_out0;
assign v$RAM$OUT_11215_out0 = v$MEM$RAM_435_out0;
assign v$BYTE$READY_13255_out0 = v$RX$BYTE$READY_2436_out0;
assign v$BYTE$RECEIVED_13441_out0 = v$RECEIVER$STREAM_564_out0;
assign v$SHIFHT$ENABLE_13500_out0 = v$G28_2098_out0;
assign v$SHIFHT$ENABLE_13501_out0 = v$G28_2099_out0;
assign v$SHIFHT$ENABLE_13502_out0 = v$G28_2100_out0;
assign v$SHIFHT$ENABLE_13503_out0 = v$G28_2101_out0;
assign v$EQ3_13504_out0 = v$Q_1153_out0 == 2'h3;
assign v$EQ3_13505_out0 = v$Q_1154_out0 == 2'h3;
assign v$DIV$INSTRUCTION_13635_out0 = v$DIV$INSTRUCTION_11296_out0;
assign v$DIV$INSTRUCTION_13636_out0 = v$DIV$INSTRUCTION_11297_out0;
assign v$EQ6_19_out0 = v$4BITCOUNTER_317_out0 == 2'h2;
assign v$R3_74_out0 = v$R3TEST_117_out0;
assign v$R3_75_out0 = v$R3TEST_118_out0;
assign v$NORMAL_181_out0 = v$EQ1_2540_out0;
assign v$NORMAL_182_out0 = v$EQ1_2541_out0;
assign v$LS_202_out0 = v$LS_204_out0;
assign v$LS_203_out0 = v$LS_205_out0;
assign v$Q1_307_out0 = v$_5832_out1;
assign v$Q1_308_out0 = v$_5833_out1;
assign v$RX$OVERFLOW_426_out0 = v$RX$OVERFLOW_4469_out0;
assign v$EXEC1LS_430_out0 = v$EQ2_8_out0;
assign v$EXEC1LS_431_out0 = v$EQ2_9_out0;
assign v$Q0_625_out0 = v$_5832_out0;
assign v$Q0_626_out0 = v$_5833_out0;
assign v$IR_640_out0 = v$IR_1871_out0;
assign v$IR_641_out0 = v$IR_1872_out0;
assign v$G7_1197_out0 = v$G11_8652_out0 && v$G12_2270_out0;
assign v$UNUSED3_1681_out0 = v$SHIFHT$ENABLE_13503_out0;
assign v$9_1700_out0 = v$G8_10609_out0;
assign v$9_1701_out0 = v$G8_10610_out0;
assign v$9_1702_out0 = v$G8_10611_out0;
assign v$9_1703_out0 = v$G8_10612_out0;
assign v$STALL$DUAL$CORE_1739_out0 = v$STALL$DUAL$CORE_3128_out0;
assign v$EQ9_2007_out0 = v$4BITCOUNTER_320_out0 == 2'h0;
assign v$R1_2056_out0 = v$R1TEST_10498_out0;
assign v$R1_2057_out0 = v$R1TEST_10499_out0;
assign v$G5_2584_out0 = ((v$G6_1159_out0 && !v$Q_293_out0) || (!v$G6_1159_out0) && v$Q_293_out0);
assign v$G5_2585_out0 = ((v$G6_1160_out0 && !v$Q_297_out0) || (!v$G6_1160_out0) && v$Q_297_out0);
assign v$G5_2586_out0 = ((v$G6_1161_out0 && !v$Q_301_out0) || (!v$G6_1161_out0) && v$Q_301_out0);
assign v$G5_2587_out0 = ((v$G6_1162_out0 && !v$Q_305_out0) || (!v$G6_1162_out0) && v$Q_305_out0);
assign v$R0_2850_out0 = v$R0TEST_7005_out0;
assign v$R0_2851_out0 = v$R0TEST_7006_out0;
assign v$G1_2911_out0 = v$EQ4_1142_out0 && v$G2_10278_out0;
assign v$EN_2919_out0 = v$EN_10451_out0;
assign v$EN_2920_out0 = v$EN_10451_out0;
assign v$EN_2921_out0 = v$EN_10451_out0;
assign v$EN_2922_out0 = v$EN_10451_out0;
assign v$EN_2923_out0 = v$EN_10452_out0;
assign v$EN_2924_out0 = v$EN_10452_out0;
assign v$EN_2925_out0 = v$EN_10452_out0;
assign v$EN_2926_out0 = v$EN_10452_out0;
assign v$EN_2927_out0 = v$EN_10453_out0;
assign v$EN_2928_out0 = v$EN_10453_out0;
assign v$EN_2929_out0 = v$EN_10453_out0;
assign v$EN_2930_out0 = v$EN_10453_out0;
assign v$EN_2931_out0 = v$EN_10454_out0;
assign v$EN_2932_out0 = v$EN_10454_out0;
assign v$EN_2933_out0 = v$EN_10454_out0;
assign v$EN_2934_out0 = v$EN_10454_out0;
assign v$START_3027_out0 = v$EQ4_611_out0;
assign v$START_3028_out0 = v$EQ4_612_out0;
assign v$RAM$OUT_3033_out0 = v$RAM$OUT_10335_out0;
assign v$RAM$OUT_3034_out0 = v$RAM$OUT_10336_out0;
assign v$G36_3135_out0 = !(v$G38_3903_out0 || v$G37_6900_out0);
assign v$G36_3136_out0 = !(v$G38_3904_out0 || v$G37_6901_out0);
assign v$G36_3137_out0 = !(v$G38_3905_out0 || v$G37_6902_out0);
assign v$G36_3138_out0 = !(v$G38_3906_out0 || v$G37_6903_out0);
assign v$EXEC2LS_3188_out0 = v$EQ3_13504_out0;
assign v$EXEC2LS_3189_out0 = v$EQ3_13505_out0;
assign v$UNUSED1_3220_out0 = v$SHIFHT$ENABLE_13502_out0;
assign v$EQ6_3257_out0 = v$4BITCOUNTER_319_out0 == 2'h0;
assign v$STALL$DUAL$CORE_3265_out0 = v$STALL$DUAL$CORE_3128_out0;
assign v$DIV$INSTRUCTION_3296_out0 = v$DIV$INSTRUCTION_13635_out0;
assign v$DIV$INSTRUCTION_3297_out0 = v$DIV$INSTRUCTION_13636_out0;
assign v$G7_6862_out0 = v$EQ_4835_out0 && v$G8_10769_out0;
assign v$G7_6863_out0 = v$EQ_4836_out0 && v$G8_10770_out0;
assign v$D_7679_out0 = v$G3_6894_out0;
assign v$D_7683_out0 = v$G3_6895_out0;
assign v$D_7687_out0 = v$G3_6896_out0;
assign v$D_7691_out0 = v$G3_6897_out0;
assign v$SHIFT$ENABLE_8684_out0 = v$SHIFHT$ENABLE_13500_out0;
assign v$EQ2_9795_out0 = v$4BITCOUNTER_317_out0 == 2'h1;
assign v$_10287_out0 = { v$Q0_4470_out0,v$Q1_6906_out0 };
assign v$_10288_out0 = { v$Q0_4471_out0,v$Q1_6907_out0 };
assign v$_10289_out0 = { v$Q0_4472_out0,v$Q1_6908_out0 };
assign v$_10290_out0 = { v$Q0_4473_out0,v$Q1_6909_out0 };
assign v$BYTE$READY_10558_out0 = v$BYTE$READY_7021_out0;
assign v$G10_10711_out0 = v$G4_6914_out0 && v$Q1_2112_out0;
assign v$R2_10904_out0 = v$R2TEST_10987_out0;
assign v$R2_10905_out0 = v$R2TEST_10988_out0;
assign v$EQ2_10981_out0 = v$4BITCOUNTER_318_out0 == 2'h0;
assign v$RESET_11174_out0 = v$G8_10609_out0;
assign v$RESET_11175_out0 = v$G8_10609_out0;
assign v$RESET_11176_out0 = v$G8_10609_out0;
assign v$RESET_11177_out0 = v$G8_10609_out0;
assign v$RESET_11178_out0 = v$G8_10610_out0;
assign v$RESET_11179_out0 = v$G8_10610_out0;
assign v$RESET_11180_out0 = v$G8_10610_out0;
assign v$RESET_11181_out0 = v$G8_10610_out0;
assign v$RESET_11182_out0 = v$G8_10611_out0;
assign v$RESET_11183_out0 = v$G8_10611_out0;
assign v$RESET_11184_out0 = v$G8_10611_out0;
assign v$RESET_11185_out0 = v$G8_10611_out0;
assign v$RESET_11186_out0 = v$G8_10612_out0;
assign v$RESET_11187_out0 = v$G8_10612_out0;
assign v$RESET_11188_out0 = v$G8_10612_out0;
assign v$RESET_11189_out0 = v$G8_10612_out0;
assign v$G9_13655_out0 = v$G6_4818_out0 && v$_2983_out1;
assign v$BYTE$RECEIVED_13796_out0 = v$BYTE$RECEIVED_13441_out0;
assign v$FLOATING$INS_13797_out0 = v$FLOATING$INSTRUCTION_10391_out0;
assign v$FLOATING$INS_13798_out0 = v$FLOATING$INSTRUCTION_10392_out0;
assign v$R3_33_out0 = v$R3_74_out0;
assign v$R3_34_out0 = v$R3_75_out0;
assign v$MUX1_650_out0 = v$G1_2911_out0 ? v$C4_10619_out0 : v$FF2_11062_out0;
assign v$G1_1167_out0 = ! v$Q0_625_out0;
assign v$G1_1168_out0 = ! v$Q0_626_out0;
assign v$FLAOTING$INSTRUCTION_1859_out0 = v$FLOATING$INS_13797_out0;
assign v$FLAOTING$INSTRUCTION_1860_out0 = v$FLOATING$INS_13798_out0;
assign v$STALL$DUAL$CORE_1959_out0 = v$STALL$DUAL$CORE_1739_out0;
assign v$BYTE$RECEIVED_2231_out0 = v$BYTE$RECEIVED_13796_out0;
assign v$R0_2537_out0 = v$R0_2850_out0;
assign v$R0_2538_out0 = v$R0_2851_out0;
assign v$RAM$OUT_2628_out0 = v$RAM$OUT_3033_out0;
assign v$RAM$OUT_2629_out0 = v$RAM$OUT_3034_out0;
assign v$R1_2630_out0 = v$R1_2056_out0;
assign v$R1_2631_out0 = v$R1_2057_out0;
assign v$G1_2700_out0 = v$RESET_11174_out0 && v$D_7679_out0;
assign v$G1_2701_out0 = v$RESET_11175_out0 && v$D_7680_out0;
assign v$G1_2703_out0 = v$RESET_11177_out0 && v$D_7682_out0;
assign v$G1_2704_out0 = v$RESET_11178_out0 && v$D_7683_out0;
assign v$G1_2705_out0 = v$RESET_11179_out0 && v$D_7684_out0;
assign v$G1_2707_out0 = v$RESET_11181_out0 && v$D_7686_out0;
assign v$G1_2708_out0 = v$RESET_11182_out0 && v$D_7687_out0;
assign v$G1_2709_out0 = v$RESET_11183_out0 && v$D_7688_out0;
assign v$G1_2711_out0 = v$RESET_11185_out0 && v$D_7690_out0;
assign v$G1_2712_out0 = v$RESET_11186_out0 && v$D_7691_out0;
assign v$G1_2713_out0 = v$RESET_11187_out0 && v$D_7692_out0;
assign v$G1_2715_out0 = v$RESET_11189_out0 && v$D_7694_out0;
assign v$BYTE$READY_2852_out0 = v$BYTE$READY_10558_out0;
assign v$LS_2864_out0 = v$LS_202_out0;
assign v$LS_2865_out0 = v$LS_203_out0;
assign v$IR_2901_out0 = v$IR_640_out0;
assign v$IR_2902_out0 = v$IR_641_out0;
assign v$_2960_out0 = { v$_10287_out0,v$Q2_6880_out0 };
assign v$_2961_out0 = { v$_10288_out0,v$Q2_6881_out0 };
assign v$_2962_out0 = { v$_10289_out0,v$Q2_6882_out0 };
assign v$_2963_out0 = { v$_10290_out0,v$Q2_6883_out0 };
assign v$G6_4531_out0 = v$G10_10711_out0 || v$G3_3343_out0;
assign v$DIV$INSTRUCTION_4614_out0 = v$DIV$INSTRUCTION_3296_out0;
assign v$DIV$INSTRUCTION_4615_out0 = v$DIV$INSTRUCTION_3297_out0;
assign v$STALL$DUAL$CORE_4696_out0 = v$STALL$DUAL$CORE_1739_out0;
assign v$G2_6791_out0 = ! v$Q1_307_out0;
assign v$G2_6792_out0 = ! v$Q1_308_out0;
assign v$EXEC1LS_6795_out0 = v$EXEC1LS_430_out0;
assign v$EXEC1LS_6796_out0 = v$EXEC1LS_431_out0;
assign v$G13_7083_out0 = v$Q0_625_out0 && v$Q1_307_out0;
assign v$G13_7084_out0 = v$Q0_626_out0 && v$Q1_308_out0;
assign v$D_7681_out0 = v$G5_2584_out0;
assign v$D_7685_out0 = v$G5_2585_out0;
assign v$D_7689_out0 = v$G5_2586_out0;
assign v$D_7693_out0 = v$G5_2587_out0;
assign v$IR_7706_out0 = v$IR_640_out0;
assign v$IR_7707_out0 = v$IR_641_out0;
assign v$R2_10556_out0 = v$R2_10904_out0;
assign v$R2_10557_out0 = v$R2_10905_out0;
assign v$EXEC2LS_10979_out0 = v$EXEC2LS_3188_out0;
assign v$EXEC2LS_10980_out0 = v$EXEC2LS_3189_out0;
assign v$STALL$DUAL$CORE_12235_out0 = v$STALL$DUAL$CORE_3265_out0;
assign v$G9_13340_out0 = v$G7_6862_out0 && v$EXEC1LS_430_out0;
assign v$G9_13341_out0 = v$G7_6863_out0 && v$EXEC1LS_431_out0;
assign v$START_13394_out0 = v$START_3027_out0;
assign v$START_13395_out0 = v$START_3028_out0;
assign v$NORMAL_13429_out0 = v$NORMAL_181_out0;
assign v$NORMAL_13430_out0 = v$NORMAL_182_out0;
assign v$9_13623_out0 = v$9_1700_out0;
assign v$9_13624_out0 = v$9_1701_out0;
assign v$9_13625_out0 = v$9_1702_out0;
assign v$9_13626_out0 = v$9_1703_out0;
assign v$_4_out0 = v$IR_2901_out0[14:12];
assign v$_5_out0 = v$IR_2902_out0[14:12];
assign v$R3_27_out0 = v$R3_33_out0;
assign v$R3_28_out0 = v$R3_34_out0;
assign v$UNUSED_123_out0 = v$9_13625_out0;
assign v$G9_223_out0 = v$G6_4531_out0 || v$G7_1197_out0;
assign v$START_392_out0 = v$START_13394_out0;
assign v$START_393_out0 = v$START_13395_out0;
assign v$9_417_out0 = v$9_13624_out0;
assign v$LS_1202_out0 = v$LS_2864_out0;
assign v$LS_1203_out0 = v$LS_2865_out0;
assign v$G7_1684_out0 = v$G1_1167_out0 && v$Q1_307_out0;
assign v$G7_1685_out0 = v$G1_1168_out0 && v$Q1_308_out0;
assign v$G3_1720_out0 = ! v$FLAOTING$INSTRUCTION_1859_out0;
assign v$G3_1721_out0 = ! v$FLAOTING$INSTRUCTION_1860_out0;
assign v$R2_1726_out0 = v$R2_10556_out0;
assign v$R2_1727_out0 = v$R2_10557_out0;
assign v$RAM$OUT_1751_out0 = v$RAM$OUT_2628_out0;
assign v$RAM$OUT_1752_out0 = v$RAM$OUT_2629_out0;
assign v$UNUSED2_2424_out0 = v$9_13626_out0;
assign v$_2599_out0 = v$IR_2901_out0[1:0];
assign v$_2600_out0 = v$IR_2902_out0[1:0];
assign v$G1_2702_out0 = v$RESET_11176_out0 && v$D_7681_out0;
assign v$G1_2706_out0 = v$RESET_11180_out0 && v$D_7685_out0;
assign v$G1_2710_out0 = v$RESET_11184_out0 && v$D_7689_out0;
assign v$G1_2714_out0 = v$RESET_11188_out0 && v$D_7693_out0;
assign v$R1_2723_out0 = v$R1_2630_out0;
assign v$R1_2724_out0 = v$R1_2631_out0;
assign v$_2773_out0 = { v$_2960_out0,v$Q3_10518_out0 };
assign v$_2774_out0 = { v$_2961_out0,v$Q3_10519_out0 };
assign v$_2775_out0 = { v$_2962_out0,v$Q3_10520_out0 };
assign v$_2776_out0 = { v$_2963_out0,v$Q3_10521_out0 };
assign v$G2_3221_out0 = ! v$9_13623_out0;
assign v$EXEC2LS_3231_out0 = v$EXEC2LS_10979_out0;
assign v$EXEC2LS_3232_out0 = v$EXEC2LS_10980_out0;
assign v$wen$ram_4595_out0 = v$G9_13340_out0;
assign v$wen$ram_4596_out0 = v$G9_13341_out0;
assign v$IR1_6873_out0 = v$IR_7706_out0;
assign v$BIT_6918_out0 = v$MUX1_650_out0;
assign v$EXEC1_7029_out0 = v$EXEC1LS_6795_out0;
assign v$EXEC1_7030_out0 = v$EXEC1LS_6796_out0;
assign v$_7095_out0 = v$IR_2901_out0[15:15];
assign v$_7096_out0 = v$IR_2902_out0[15:15];
assign v$STALL$dual$core_8742_out0 = v$STALL$DUAL$CORE_1959_out0;
assign v$BYTE$RECEIVED_8819_out0 = v$BYTE$RECEIVED_2231_out0;
assign v$BYTE$RECEIVED_8820_out0 = v$BYTE$RECEIVED_2231_out0;
assign v$NORMAL_10256_out0 = v$NORMAL_13429_out0;
assign v$NORMAL_10257_out0 = v$NORMAL_13430_out0;
assign v$_10371_out0 = { v$STALL$DUAL$CORE_4696_out0,v$C_1808_out0 };
assign v$EXEC1LS_10506_out0 = v$EXEC1LS_6795_out0;
assign v$EXEC1LS_10507_out0 = v$EXEC1LS_6796_out0;
assign v$_10791_out0 = v$IR_2901_out0[11:10];
assign v$_10792_out0 = v$IR_2902_out0[11:10];
assign v$G5_10914_out0 = v$Q0_625_out0 && v$G2_6791_out0;
assign v$G5_10915_out0 = v$Q0_626_out0 && v$G2_6792_out0;
assign v$BYTE$RECEIVED_11192_out0 = v$BYTE$RECEIVED_2231_out0;
assign v$STORE_12245_out0 = v$G9_13340_out0;
assign v$STORE_12246_out0 = v$G9_13341_out0;
assign v$R0_13295_out0 = v$R0_2537_out0;
assign v$R0_13296_out0 = v$R0_2538_out0;
assign v$IR0_13305_out0 = v$IR_7707_out0;
assign v$IR_13480_out0 = v$IR_2901_out0;
assign v$IR_13481_out0 = v$IR_2902_out0;
assign v$G3_13641_out0 = v$G1_1167_out0 && v$G2_6791_out0;
assign v$G3_13642_out0 = v$G1_1168_out0 && v$G2_6792_out0;
assign v$IR_105_out0 = v$IR_13480_out0;
assign v$IR_106_out0 = v$IR_13481_out0;
assign v$_224_out0 = v$RAM$OUT_1751_out0[11:0];
assign v$_224_out1 = v$RAM$OUT_1751_out0[15:4];
assign v$_225_out0 = v$RAM$OUT_1752_out0[11:0];
assign v$_225_out1 = v$RAM$OUT_1752_out0[15:4];
assign v$G1_277_out0 = v$EQ2_9795_out0 && v$G2_3221_out0;
assign v$R13_375_out0 = v$R3_27_out0;
assign v$R11_398_out0 = v$R1_2723_out0;
assign v$_533_out0 = { v$G1_10810_out0,v$G9_223_out0 };
assign v$OP_621_out0 = v$_4_out0;
assign v$OP_622_out0 = v$_5_out0;
assign v$D_2108_out0 = v$_10791_out0;
assign v$D_2109_out0 = v$_10792_out0;
assign v$G16_2310_out0 = ! v$STORE_12245_out0;
assign v$G16_2311_out0 = ! v$STORE_12246_out0;
assign v$_2422_out0 = v$IR_13480_out0[8:8];
assign v$_2423_out0 = v$IR_13481_out0[8:8];
assign v$IR15_2464_out0 = v$_7095_out0;
assign v$IR15_2465_out0 = v$_7096_out0;
assign v$G8_2644_out0 = ! v$9_417_out0;
assign v$_2846_out0 = v$IR_13480_out0[4:0];
assign v$_2847_out0 = v$IR_13481_out0[4:0];
assign v$G6_2905_out0 = v$G3_13641_out0 || v$G7_1684_out0;
assign v$G6_2906_out0 = v$G3_13642_out0 || v$G7_1685_out0;
assign v$LS1_3169_out0 = v$LS_1202_out0;
assign v$BIT$IN1_3209_out0 = v$BIT_6918_out0;
assign v$NORMAL_3353_out0 = v$NORMAL_10256_out0;
assign v$NORMAL_3354_out0 = v$NORMAL_10257_out0;
assign v$R00_3807_out0 = v$R0_13296_out0;
assign v$_3942_out0 = v$IR_13480_out0[7:4];
assign v$_3943_out0 = v$IR_13481_out0[7:4];
assign v$LS0_4548_out0 = v$LS_1203_out0;
assign v$_4837_out0 = v$IR_13480_out0[9:9];
assign v$_4838_out0 = v$IR_13481_out0[9:9];
assign v$SEL1_5798_out0 = v$IR_13480_out0[15:12];
assign v$SEL1_5799_out0 = v$IR_13481_out0[15:12];
assign v$R02_6966_out0 = v$R2_1727_out0;
assign v$WEN$RAM_7079_out0 = v$wen$ram_4595_out0;
assign v$WEN$RAM_7080_out0 = v$wen$ram_4596_out0;
assign v$EN_7094_out0 = v$STALL$dual$core_8742_out0;
assign v$BYTE$RECEIVED_7101_out0 = v$BYTE$RECEIVED_8819_out0;
assign v$BYTE$RECEIVED_7102_out0 = v$BYTE$RECEIVED_8820_out0;
assign v$M_7177_out0 = v$_2599_out0;
assign v$M_7178_out0 = v$_2600_out0;
assign v$R12_10714_out0 = v$R2_1726_out0;
assign v$EXEC1_10763_out0 = v$EXEC1_7029_out0;
assign v$EXEC1_10764_out0 = v$EXEC1_7030_out0;
assign v$A_10822_out0 = v$_10371_out0;
assign v$EXEC1LS_10843_out0 = v$EXEC1LS_10506_out0;
assign v$EXEC1LS_10844_out0 = v$EXEC1LS_10507_out0;
assign v$_11163_out0 = v$IR_13480_out0[3:2];
assign v$_11164_out0 = v$IR_13481_out0[3:2];
assign v$R10_11216_out0 = v$R0_13295_out0;
assign v$8BITCOUNTER_13281_out0 = v$_2773_out0;
assign v$8BITCOUNTER_13282_out0 = v$_2774_out0;
assign v$8BITCOUNTER_13283_out0 = v$_2775_out0;
assign v$8BITCOUNTER_13284_out0 = v$_2776_out0;
assign v$R03_13304_out0 = v$R3_28_out0;
assign v$EXEC2LS_13558_out0 = v$EXEC2LS_3231_out0;
assign v$EXEC2LS_13559_out0 = v$EXEC2LS_3232_out0;
assign v$WRITE$EN_13653_out0 = v$wen$ram_4595_out0;
assign v$WRITE$EN_13654_out0 = v$wen$ram_4596_out0;
assign v$R01_13752_out0 = v$R1_2724_out0;
assign v$_61_out0 = v$A_10822_out0[10:10];
assign v$_172_out0 = v$A_10822_out0[7:7];
assign v$_180_out0 = v$A_10822_out0[3:3];
assign v$B_273_out0 = v$_3942_out0;
assign v$B_274_out0 = v$_3943_out0;
assign v$_288_out0 = v$A_10822_out0[2:2];
assign v$EQ1_315_out0 = v$_224_out1 == 4'h0;
assign v$EQ1_316_out0 = v$_225_out1 == 4'h0;
assign v$G15_1855_out0 = !(v$EXEC1_10763_out0 || v$FF1_48_out0);
assign v$G15_1856_out0 = !(v$EXEC1_10764_out0 || v$FF1_49_out0);
assign v$EQ1_1857_out0 = v$SEL1_5798_out0 == 4'h1;
assign v$EQ1_1858_out0 = v$SEL1_5799_out0 == 4'h1;
assign v$_1876_out0 = v$A_10822_out0[11:11];
assign v$EQ6_1966_out0 = v$_224_out1 == 4'h5;
assign v$EQ6_1967_out0 = v$_225_out1 == 4'h5;
assign v$_2023_out0 = v$A_10822_out0[5:5];
assign v$EXEC2_2110_out0 = v$EXEC2LS_13558_out0;
assign v$EXEC2_2111_out0 = v$EXEC2LS_13559_out0;
assign v$EQ4_2149_out0 = v$8BITCOUNTER_13281_out0 == 4'h0;
assign v$_2269_out0 = v$A_10822_out0[8:8];
assign v$EQ9_2390_out0 = v$_224_out1 == 4'h3;
assign v$EQ9_2391_out0 = v$_225_out1 == 4'h3;
assign v$EQ8_2453_out0 = v$_224_out1 == 4'h7;
assign v$EQ8_2454_out0 = v$_225_out1 == 4'h7;
assign v$EQ11_2456_out0 = v$_224_out1 == 4'h1;
assign v$EQ11_2457_out0 = v$_225_out1 == 4'h1;
assign v$IN_2466_out0 = v$BIT$IN1_3209_out0;
assign v$ADRESS_2542_out0 = v$_224_out0;
assign v$ADRESS_2543_out0 = v$_225_out0;
assign v$G21_2656_out0 = ! v$WEN$RAM_7079_out0;
assign v$G21_2657_out0 = ! v$WEN$RAM_7080_out0;
assign v$WEN_2765_out0 = v$WRITE$EN_13653_out0;
assign v$WEN_2766_out0 = v$WRITE$EN_13654_out0;
assign v$EXEC2LS_2844_out0 = v$EXEC2LS_13558_out0;
assign v$EXEC2LS_2845_out0 = v$EXEC2LS_13559_out0;
assign v$EQ8_2874_out0 = v$8BITCOUNTER_13284_out0 == 4'h0;
assign v$SEL1_2914_out0 = v$_224_out0[9:9];
assign v$SEL1_2915_out0 = v$_225_out0[9:9];
assign v$EQ3_2966_out0 = v$SEL1_5798_out0 == 4'h9;
assign v$EQ3_2967_out0 = v$SEL1_5799_out0 == 4'h9;
assign v$_3124_out0 = v$A_10822_out0[1:1];
assign v$EXEC2_3170_out0 = v$NORMAL_3353_out0;
assign v$EXEC2_3171_out0 = v$NORMAL_3354_out0;
assign v$EQ4_3227_out0 = v$SEL1_5798_out0 == 4'h8;
assign v$EQ4_3228_out0 = v$SEL1_5799_out0 == 4'h8;
assign v$_3271_out0 = v$A_10822_out0[4:4];
assign v$EQ7_3307_out0 = v$_224_out1 == 4'h6;
assign v$EQ7_3308_out0 = v$_225_out1 == 4'h6;
assign v$exec1ls_3341_out0 = v$EXEC1LS_10843_out0;
assign v$exec1ls_3342_out0 = v$EXEC1LS_10844_out0;
assign v$EXEC1LS_4697_out0 = v$EXEC1LS_10843_out0;
assign v$EXEC1LS_4698_out0 = v$EXEC1LS_10844_out0;
assign v$EQ5_4860_out0 = v$_224_out1 == 4'h4;
assign v$EQ5_4861_out0 = v$_225_out1 == 4'h4;
assign v$K_5792_out0 = v$_2846_out0;
assign v$K_5793_out0 = v$_2847_out0;
assign v$_7081_out0 = { v$BYTE$RECEIVED_7101_out0,v$C1_13277_out0 };
assign v$_7082_out0 = { v$BYTE$RECEIVED_7102_out0,v$C1_13278_out0 };
assign v$NORMAL_7114_out0 = v$NORMAL_3353_out0;
assign v$NORMAL_7115_out0 = v$NORMAL_3354_out0;
assign v$EXEC1_7128_out0 = v$EXEC1LS_10843_out0;
assign v$EXEC1_7129_out0 = v$EXEC1LS_10844_out0;
assign v$EQ3_7145_out0 = v$_224_out1 == 4'h2;
assign v$EQ3_7146_out0 = v$_225_out1 == 4'h2;
assign v$C_8653_out0 = v$_4837_out0;
assign v$C_8654_out0 = v$_4838_out0;
assign v$SHIFT_8661_out0 = v$_11163_out0;
assign v$SHIFT_8662_out0 = v$_11164_out0;
assign v$D_8752_out0 = v$D_2108_out0;
assign v$D_8753_out0 = v$D_2109_out0;
assign v$_9791_out0 = { v$C1_13277_out0,v$BYTE$RECEIVED_7101_out0 };
assign v$_9792_out0 = { v$C1_13278_out0,v$BYTE$RECEIVED_7102_out0 };
assign v$EQ1_10329_out0 = v$8BITCOUNTER_13282_out0 == 4'h0;
assign v$LDR$STR0_10349_out0 = v$LS0_4548_out0;
assign v$AD2_10699_out0 = v$M_7177_out0;
assign v$AD2_10700_out0 = v$M_7178_out0;
assign v$IR_10816_out0 = v$IR_105_out0;
assign v$IR_10817_out0 = v$IR_106_out0;
assign v$OP_11223_out0 = v$OP_621_out0;
assign v$OP_11224_out0 = v$OP_622_out0;
assign v$_11243_out0 = v$A_10822_out0[9:9];
assign v$S_11300_out0 = v$_2422_out0;
assign v$S_11301_out0 = v$_2423_out0;
assign v$_13397_out0 = v$A_10822_out0[6:6];
assign v$_13563_out0 = v$A_10822_out0[0:0];
assign v$LDR$STR1_13616_out0 = v$LS1_3169_out0;
assign v$EQ7_13769_out0 = v$8BITCOUNTER_13283_out0 == 4'h0;
assign v$AD1_13774_out0 = v$D_2108_out0;
assign v$AD1_13775_out0 = v$D_2109_out0;
assign v$BIT$STREAM$IN_13_out0 = v$IN_2466_out0;
assign v$G4_381_out0 = v$EQ3_2966_out0 || v$EQ4_3227_out0;
assign v$G4_382_out0 = v$EQ3_2967_out0 || v$EQ4_3228_out0;
assign v$G20_598_out0 = v$EXEC1_10763_out0 && v$G21_2656_out0;
assign v$G20_599_out0 = v$EXEC1_10764_out0 && v$G21_2657_out0;
assign v$EXEC20_629_out0 = v$EXEC2_2111_out0;
assign v$B_1155_out0 = v$B_273_out0;
assign v$B_1156_out0 = v$B_274_out0;
assign v$EQ6_1686_out0 = v$OP_11223_out0 == 3'h5;
assign v$EQ6_1687_out0 = v$OP_11224_out0 == 3'h5;
assign v$_1724_out0 = v$IR_10816_out0[14:14];
assign v$_1725_out0 = v$IR_10817_out0[14:14];
assign v$JMI_1939_out0 = v$EQ6_1966_out0;
assign v$JMI_1940_out0 = v$EQ6_1967_out0;
assign v$EXEC2_2010_out0 = v$EXEC2_3170_out0;
assign v$EXEC2_2011_out0 = v$EXEC2_3171_out0;
assign v$NORMAL0_2307_out0 = v$NORMAL_7115_out0;
assign v$EXEC10_2329_out0 = v$exec1ls_3342_out0;
assign v$ADRESS_2339_out0 = v$ADRESS_2542_out0;
assign v$ADRESS_2340_out0 = v$ADRESS_2543_out0;
assign v$_2430_out0 = v$IR_10816_out0[15:15];
assign v$_2431_out0 = v$IR_10817_out0[15:15];
assign v$_2470_out0 = v$IR_10816_out0[13:13];
assign v$_2471_out0 = v$IR_10817_out0[13:13];
assign v$K_2636_out0 = v$K_5792_out0;
assign v$K_2637_out0 = v$K_5793_out0;
assign v$G2_2652_out0 = v$EQ9_2390_out0 || v$EQ10_2320_out0;
assign v$G2_2653_out0 = v$EQ9_2391_out0 || v$EQ10_2321_out0;
assign v$SUB_2695_out0 = v$EQ3_2966_out0;
assign v$SUB_2696_out0 = v$EQ3_2967_out0;
assign v$G5_2756_out0 = ! v$SEL1_2914_out0;
assign v$G5_2757_out0 = ! v$SEL1_2915_out0;
assign v$_2831_out0 = v$AD2_10699_out0[0:0];
assign v$_2831_out1 = v$AD2_10699_out0[1:1];
assign v$_2832_out0 = v$AD2_10700_out0[0:0];
assign v$_2832_out1 = v$AD2_10700_out0[1:1];
assign v$_2860_out0 = v$IR_10816_out0[12:12];
assign v$_2861_out0 = v$IR_10817_out0[12:12];
assign v$EQ8_2951_out0 = v$OP_11223_out0 == 3'h7;
assign v$EQ8_2952_out0 = v$OP_11224_out0 == 3'h7;
assign v$MULTI$OPCODE_3020_out0 = v$EQ1_1857_out0;
assign v$MULTI$OPCODE_3021_out0 = v$EQ1_1858_out0;
assign v$EXEC1_3038_out0 = v$EXEC1_7128_out0;
assign v$EXEC1_3039_out0 = v$EXEC1_7129_out0;
assign v$EXEC2LS_3081_out0 = v$EXEC2LS_2844_out0;
assign v$EXEC2LS_3082_out0 = v$EXEC2LS_2845_out0;
assign v$_3897_out0 = v$IR_10816_out0[9:0];
assign v$_3897_out1 = v$IR_10816_out0[15:6];
assign v$_3898_out0 = v$IR_10817_out0[9:0];
assign v$_3898_out1 = v$IR_10817_out0[15:6];
assign v$EXEC11_4528_out0 = v$exec1ls_3341_out0;
assign v$FLOAT_4603_out0 = v$EQ3_7145_out0;
assign v$FLOAT_4604_out0 = v$EQ3_7146_out0;
assign v$G25_4658_out0 = v$EQ8_2874_out0 && v$EQ9_2007_out0;
assign v$NORMAL1_6790_out0 = v$NORMAL_7114_out0;
assign v$REN1_6874_out0 = v$LDR$STR1_13616_out0;
assign v$_6876_out0 = v$AD1_13774_out0[0:0];
assign v$_6876_out1 = v$AD1_13774_out0[1:1];
assign v$_6877_out0 = v$AD1_13775_out0[0:0];
assign v$_6877_out1 = v$AD1_13775_out0[1:1];
assign v$EQ1_7098_out0 = v$OP_11223_out0 == 3'h0;
assign v$EQ1_7099_out0 = v$OP_11224_out0 == 3'h0;
assign v$EQ3_7126_out0 = v$OP_11223_out0 == 3'h2;
assign v$EQ3_7127_out0 = v$OP_11224_out0 == 3'h2;
assign v$JMP_8825_out0 = v$EQ5_4860_out0;
assign v$JMP_8826_out0 = v$EQ5_4861_out0;
assign v$EQ4_10345_out0 = v$OP_11223_out0 == 3'h3;
assign v$EQ4_10346_out0 = v$OP_11224_out0 == 3'h3;
assign v$STP_10352_out0 = v$EQ8_2453_out0;
assign v$STP_10353_out0 = v$EQ8_2454_out0;
assign v$EQ5_10364_out0 = v$OP_11223_out0 == 3'h4;
assign v$EQ5_10365_out0 = v$OP_11224_out0 == 3'h4;
assign v$EQ7_10399_out0 = v$OP_11223_out0 == 3'h6;
assign v$EQ7_10400_out0 = v$OP_11224_out0 == 3'h6;
assign v$JEQ_10496_out0 = v$EQ7_3307_out0;
assign v$JEQ_10497_out0 = v$EQ7_3308_out0;
assign v$RD_10522_out0 = v$D_8752_out0;
assign v$RD_10523_out0 = v$D_8753_out0;
assign v$EXEC2LS_10549_out0 = v$EXEC2_2110_out0;
assign v$SHIFT_10615_out0 = v$SHIFT_8661_out0;
assign v$SHIFT_10616_out0 = v$SHIFT_8662_out0;
assign v$G22_10620_out0 = v$EQ7_13769_out0 && v$EQ6_3257_out0;
assign v$EXEC1LS_10703_out0 = v$EXEC1LS_4697_out0;
assign v$EXEC1LS_10704_out0 = v$EXEC1LS_4698_out0;
assign v$EQ2_10771_out0 = v$OP_11223_out0 == 3'h1;
assign v$EQ2_10772_out0 = v$OP_11224_out0 == 3'h1;
assign v$G5_10989_out0 = ! v$EQ4_2149_out0;
assign v$WEN_11038_out0 = v$WEN_2765_out0;
assign v$WEN_11039_out0 = v$WEN_2766_out0;
assign v$REN0_11136_out0 = v$LDR$STR0_10349_out0;
assign v$G1_11157_out0 = v$EQ1_315_out0 || v$EQ9_2390_out0;
assign v$G1_11158_out0 = v$EQ1_316_out0 || v$EQ9_2391_out0;
assign v$G9_13564_out0 = v$EQ2_10981_out0 && v$EQ1_10329_out0;
assign v$C_13767_out0 = v$C_8653_out0;
assign v$C_13768_out0 = v$C_8654_out0;
assign v$G8_16_out0 = v$G1_277_out0 && v$BIT$STREAM$IN_13_out0;
assign v$STP_52_out0 = v$STP_10352_out0;
assign v$STP_53_out0 = v$STP_10353_out0;
assign v$_124_out0 = { v$K_2636_out0,v$C1_606_out0 };
assign v$_125_out0 = { v$K_2637_out0,v$C1_607_out0 };
assign v$C_238_out0 = v$C_13767_out0;
assign v$C_239_out0 = v$C_13768_out0;
assign v$MUX4_376_out0 = v$_2831_out0 ? v$R1_8761_out0 : v$R0_1688_out0;
assign v$MUX4_377_out0 = v$_2832_out0 ? v$R1_8762_out0 : v$R0_1689_out0;
assign v$EXEC2_441_out0 = v$EXEC2_2010_out0;
assign v$EXEC2_442_out0 = v$EXEC2_2011_out0;
assign v$G4_1667_out0 = v$EQ1_315_out0 && v$G5_2756_out0;
assign v$G4_1668_out0 = v$EQ1_316_out0 && v$G5_2757_out0;
assign v$UART_1823_out0 = v$G2_2652_out0;
assign v$UART_1824_out0 = v$G2_2653_out0;
assign v$EXEC1_1863_out0 = v$EXEC1LS_10703_out0;
assign v$EXEC1_1864_out0 = v$EXEC1LS_10704_out0;
assign v$G3_1949_out0 = v$EQ11_2456_out0 || v$G1_11157_out0;
assign v$G3_1950_out0 = v$EQ11_2457_out0 || v$G1_11158_out0;
assign v$JEQ_2234_out0 = v$JEQ_10496_out0;
assign v$JEQ_2235_out0 = v$JEQ_10497_out0;
assign v$BIT_2328_out0 = v$BIT$STREAM$IN_13_out0;
assign v$G7_2455_out0 = v$G9_13564_out0 || v$G8_2644_out0;
assign v$MUX1_2532_out0 = v$_6876_out0 ? v$REG1_2314_out0 : v$REG0_10912_out0;
assign v$MUX1_2533_out0 = v$_6877_out0 ? v$REG1_2315_out0 : v$REG0_10913_out0;
assign v$WEN0_2588_out0 = v$WEN_11039_out0;
assign v$EXEC1_2634_out0 = v$EXEC1LS_10703_out0;
assign v$EXEC1_2635_out0 = v$EXEC1LS_10704_out0;
assign v$EXEC2_2647_out0 = v$EXEC2LS_3081_out0;
assign v$EXEC2_2648_out0 = v$EXEC2LS_3082_out0;
assign v$NOTUSED_2698_out0 = v$_3897_out1;
assign v$NOTUSED_2699_out0 = v$_3898_out1;
assign v$SUB$INSTRUCTION_2789_out0 = v$SUB_2695_out0;
assign v$SUB$INSTRUCTION_2790_out0 = v$SUB_2696_out0;
assign v$EXEC11_2830_out0 = v$EXEC11_4528_out0;
assign v$JMP_3233_out0 = v$JMP_8825_out0;
assign v$JMP_3234_out0 = v$JMP_8826_out0;
assign v$EXEC2_3241_out0 = v$EXEC2LS_3081_out0;
assign v$EXEC2_3242_out0 = v$EXEC2LS_3082_out0;
assign v$TST_3819_out0 = v$EQ8_2951_out0;
assign v$TST_3820_out0 = v$EQ8_2952_out0;
assign v$AND_3858_out0 = v$EQ7_10399_out0;
assign v$AND_3859_out0 = v$EQ7_10400_out0;
assign v$MULTI$INSTRUCTION_3953_out0 = v$MULTI$OPCODE_3020_out0;
assign v$MULTI$INSTRUCTION_3954_out0 = v$MULTI$OPCODE_3021_out0;
assign v$G24_3955_out0 = ! v$_2470_out0;
assign v$G24_3956_out0 = ! v$_2471_out0;
assign v$G3_3959_out0 = v$G4_381_out0 && v$FLOATING$INS_13797_out0;
assign v$G3_3960_out0 = v$G4_382_out0 && v$FLOATING$INS_13798_out0;
assign v$ADD_4455_out0 = v$EQ1_7098_out0;
assign v$ADD_4456_out0 = v$EQ1_7099_out0;
assign v$_4526_out0 = v$_3897_out0[8:0];
assign v$_4526_out1 = v$_3897_out0[9:1];
assign v$_4527_out0 = v$_3898_out0[8:0];
assign v$_4527_out1 = v$_3898_out0[9:1];
assign v$MUX2_4612_out0 = v$_6876_out0 ? v$REG3_4747_out0 : v$REG2_12251_out0;
assign v$MUX2_4613_out0 = v$_6877_out0 ? v$REG3_4748_out0 : v$REG2_12252_out0;
assign v$BIN_5853_out0 = v$B_1155_out0;
assign v$BIN_5854_out0 = v$B_1156_out0;
assign v$G28_6868_out0 = ! v$_1724_out0;
assign v$G28_6869_out0 = ! v$_1725_out0;
assign v$G25_6962_out0 = v$_2430_out0 && v$_1724_out0;
assign v$G25_6963_out0 = v$_2431_out0 && v$_1725_out0;
assign v$JUMPADRESS_6964_out0 = v$ADRESS_2339_out0;
assign v$JUMPADRESS_6965_out0 = v$ADRESS_2340_out0;
assign v$STARTBIT_6967_out0 = v$BIT$STREAM$IN_13_out0;
assign v$FLOAT_7676_out0 = v$FLOAT_4603_out0;
assign v$FLOAT_7677_out0 = v$FLOAT_4604_out0;
assign v$SUB_8663_out0 = v$EQ2_10771_out0;
assign v$SUB_8664_out0 = v$EQ2_10772_out0;
assign v$WEN1_8763_out0 = v$WEN_11038_out0;
assign v$EXEC10_8812_out0 = v$EXEC10_2329_out0;
assign v$MUX5_8840_out0 = v$_2831_out0 ? v$R3_4652_out0 : v$R2_3043_out0;
assign v$MUX5_8841_out0 = v$_2832_out0 ? v$R3_4653_out0 : v$R2_3044_out0;
assign v$MOV_10389_out0 = v$EQ5_10364_out0;
assign v$MOV_10390_out0 = v$EQ5_10365_out0;
assign v$ADC_10393_out0 = v$EQ3_7126_out0;
assign v$ADC_10394_out0 = v$EQ3_7127_out0;
assign v$G3_10462_out0 = v$G5_10989_out0 && v$EQ6_19_out0;
assign v$G21_10681_out0 = ! v$G22_10620_out0;
assign v$MULTI$OPCODE_11096_out0 = v$MULTI$OPCODE_3020_out0;
assign v$MULTI$OPCODE_11097_out0 = v$MULTI$OPCODE_3021_out0;
assign v$G2_12230_out0 = v$EXEC2_2010_out0 || v$EXEC2LS_3081_out0;
assign v$G2_12231_out0 = v$EXEC2_2011_out0 || v$EXEC2LS_3082_out0;
assign v$JMI_13349_out0 = v$JMI_1939_out0;
assign v$JMI_13350_out0 = v$JMI_1940_out0;
assign v$SBC_13605_out0 = v$EQ4_10345_out0;
assign v$SBC_13606_out0 = v$EQ4_10346_out0;
assign v$CMP_13609_out0 = v$EQ6_1686_out0;
assign v$CMP_13610_out0 = v$EQ6_1687_out0;
assign v$EXEC1_20_out0 = v$EXEC1_1863_out0;
assign v$EXEC1_21_out0 = v$EXEC1_1864_out0;
assign v$JMI_88_out0 = v$JMI_13349_out0;
assign v$JMI_89_out0 = v$JMI_13350_out0;
assign v$MOV_196_out0 = v$MOV_10389_out0;
assign v$MOV_197_out0 = v$MOV_10390_out0;
assign v$MUX3_313_out0 = v$_6876_out1 ? v$MUX2_4612_out0 : v$MUX1_2532_out0;
assign v$MUX3_314_out0 = v$_6877_out1 ? v$MUX2_4613_out0 : v$MUX1_2533_out0;
assign v$C_379_out0 = v$C_238_out0;
assign v$C_380_out0 = v$C_239_out0;
assign v$STALL_427_out0 = v$G3_1949_out0;
assign v$STALL_428_out0 = v$G3_1950_out0;
assign v$MUX1_534_out0 = v$C_238_out0 ? v$ROR_66_out0 : v$SHIFT_10615_out0;
assign v$MUX1_535_out0 = v$C_239_out0 ? v$ROR_67_out0 : v$SHIFT_10616_out0;
assign v$JMP_546_out0 = v$JMP_3233_out0;
assign v$JMP_547_out0 = v$JMP_3234_out0;
assign v$G18_567_out0 = v$EXEC11_2830_out0 && v$REN1_6874_out0;
assign v$FLOATING$EN$ALU_634_out0 = v$G3_3959_out0;
assign v$FLOATING$EN$ALU_635_out0 = v$G3_3960_out0;
assign v$MUX2_1145_out0 = v$G2_12230_out0 ? v$D_2108_out0 : v$M_7177_out0;
assign v$MUX2_1146_out0 = v$G2_12231_out0 ? v$D_2109_out0 : v$M_7178_out0;
assign v$EQ1_1157_out0 = v$_4526_out1 == 1'h0;
assign v$EQ1_1158_out0 = v$_4527_out1 == 1'h0;
assign v$G1_2225_out0 = ! v$TST_3819_out0;
assign v$G1_2226_out0 = ! v$TST_3820_out0;
assign v$MUX6_2341_out0 = v$_2831_out1 ? v$MUX5_8840_out0 : v$MUX4_376_out0;
assign v$MUX6_2342_out0 = v$_2832_out1 ? v$MUX5_8841_out0 : v$MUX4_377_out0;
assign v$WEN0_2646_out0 = v$WEN0_2588_out0;
assign v$G23_2840_out0 = v$G25_6962_out0 && v$G24_3955_out0;
assign v$G23_2841_out0 = v$G25_6963_out0 && v$G24_3956_out0;
assign v$G2_2891_out0 = v$EXEC1_2634_out0 && v$G3_1720_out0;
assign v$G2_2892_out0 = v$EXEC1_2635_out0 && v$G3_1721_out0;
assign v$G3_2941_out0 = v$FLOAT_7676_out0 && v$NORMAL_13429_out0;
assign v$G3_2942_out0 = v$FLOAT_7677_out0 && v$NORMAL_13430_out0;
assign v$SUB_2957_out0 = v$SUB_8663_out0;
assign v$SUB_2958_out0 = v$SUB_8664_out0;
assign v$G16_3024_out0 = v$EXEC10_8812_out0 && v$REN0_11136_out0;
assign v$_3040_out0 = { v$_2959_out1,v$BIT_2328_out0 };
assign v$JMI_3212_out0 = v$JMI_13349_out0;
assign v$JMI_3213_out0 = v$JMI_13350_out0;
assign v$CMP_3805_out0 = v$CMP_13609_out0;
assign v$CMP_3806_out0 = v$CMP_13610_out0;
assign v$JEQ_4445_out0 = v$JEQ_2234_out0;
assign v$JEQ_4446_out0 = v$JEQ_2235_out0;
assign v$JUMPADRESS_4745_out0 = v$JUMPADRESS_6964_out0;
assign v$JUMPADRESS_4746_out0 = v$JUMPADRESS_6965_out0;
assign v$SBC_4825_out0 = v$SBC_13605_out0;
assign v$SBC_4826_out0 = v$SBC_13606_out0;
assign v$G2_6884_out0 = v$S_11300_out0 && v$EXEC2_441_out0;
assign v$G2_6885_out0 = v$S_11301_out0 && v$EXEC2_442_out0;
assign v$JMP_7077_out0 = v$JMP_3233_out0;
assign v$JMP_7078_out0 = v$JMP_3234_out0;
assign v$EQ2_7091_out0 = v$_4526_out1 == 1'h1;
assign v$EQ2_7092_out0 = v$_4527_out1 == 1'h1;
assign v$EXEC2_7181_out0 = v$EXEC2_2647_out0;
assign v$EXEC2_7182_out0 = v$EXEC2_2648_out0;
assign v$TST_8735_out0 = v$TST_3819_out0;
assign v$TST_8736_out0 = v$TST_3820_out0;
assign v$JEQ_8806_out0 = v$JEQ_2234_out0;
assign v$JEQ_8807_out0 = v$JEQ_2235_out0;
assign v$G27_9793_out0 = v$_2430_out0 && v$G28_6868_out0;
assign v$G27_9794_out0 = v$_2431_out0 && v$G28_6869_out0;
assign v$Wen1_10312_out0 = v$WEN1_8763_out0;
assign v$G7_10332_out0 = v$9_13623_out0 && v$G3_10462_out0;
assign v$G35_10360_out0 = v$STARTBIT_6967_out0 && v$G36_3135_out0;
assign v$G5_10441_out0 = ! v$CMP_13609_out0;
assign v$G5_10442_out0 = ! v$CMP_13610_out0;
assign v$STP_10467_out0 = v$STP_52_out0;
assign v$STP_10468_out0 = v$STP_53_out0;
assign v$MULTI$OPCODE_10797_out0 = v$MULTI$OPCODE_11096_out0;
assign v$MULTI$OPCODE_10798_out0 = v$MULTI$OPCODE_11097_out0;
assign v$UART_10825_out0 = v$UART_1823_out0;
assign v$UART_10826_out0 = v$UART_1824_out0;
assign v$_10868_out0 = v$_4526_out0[7:0];
assign v$_10868_out1 = v$_4526_out0[8:1];
assign v$_10869_out0 = v$_4527_out0[7:0];
assign v$_10869_out1 = v$_4527_out0[8:1];
assign v$STP_10977_out0 = v$STP_52_out0;
assign v$STP_10978_out0 = v$STP_53_out0;
assign v$G6_11143_out0 = v$G4_1667_out0 && v$NORMAL_181_out0;
assign v$G6_11144_out0 = v$G4_1668_out0 && v$NORMAL_182_out0;
assign v$ADD_11193_out0 = v$ADD_4455_out0;
assign v$ADD_11194_out0 = v$ADD_4456_out0;
assign v$SUB$INSTRUCTION_11195_out0 = v$SUB$INSTRUCTION_2789_out0;
assign v$SUB$INSTRUCTION_11196_out0 = v$SUB$INSTRUCTION_2790_out0;
assign v$BYTERECEIVED_11197_out0 = v$G8_16_out0;
assign v$_13253_out0 = v$BIN_5853_out0[3:1];
assign v$_13254_out0 = v$BIN_5854_out0[3:1];
assign v$MULTI$INSTRUCTION_13323_out0 = v$MULTI$INSTRUCTION_3953_out0;
assign v$MULTI$INSTRUCTION_13324_out0 = v$MULTI$INSTRUCTION_3954_out0;
assign v$KEXTEND_13329_out0 = v$_124_out0;
assign v$KEXTEND_13330_out0 = v$_125_out0;
assign v$AND_13556_out0 = v$AND_3858_out0;
assign v$AND_13557_out0 = v$AND_3859_out0;
assign v$ADC_13614_out0 = v$ADC_10393_out0;
assign v$ADC_13615_out0 = v$ADC_10394_out0;
assign v$G3_17_out0 = v$G1_2225_out0 && v$EXEC2_441_out0;
assign v$G3_18_out0 = v$G1_2226_out0 && v$EXEC2_442_out0;
assign v$SR_371_out0 = v$MUX1_534_out0;
assign v$SR_372_out0 = v$MUX1_535_out0;
assign v$TST_409_out0 = v$TST_8735_out0;
assign v$TST_410_out0 = v$TST_8736_out0;
assign v$SR_542_out0 = v$MUX1_534_out0;
assign v$SR_543_out0 = v$MUX1_535_out0;
assign v$MULTI$INSTRUCTION_619_out0 = v$MULTI$INSTRUCTION_13323_out0;
assign v$MULTI$INSTRUCTION_620_out0 = v$MULTI$INSTRUCTION_13324_out0;
assign v$STORE_1195_out0 = v$EQ1_1157_out0;
assign v$STORE_1196_out0 = v$EQ1_1158_out0;
assign v$DOUT1_1207_out0 = v$MUX3_313_out0;
assign v$DOUT1_1208_out0 = v$MUX3_314_out0;
assign v$DOUT2_1733_out0 = v$MUX6_2341_out0;
assign v$DOUT2_1734_out0 = v$MUX6_2342_out0;
assign v$ENABLE_1757_out0 = v$G7_10332_out0;
assign v$STALL_1758_out0 = v$STALL_427_out0;
assign v$STALL_1759_out0 = v$STALL_428_out0;
assign v$ADC_1821_out0 = v$ADC_13614_out0;
assign v$ADC_1822_out0 = v$ADC_13615_out0;
assign v$SR_1956_out0 = v$MUX1_534_out0;
assign v$SR_1957_out0 = v$MUX1_535_out0;
assign v$ENABLE_2018_out0 = v$G35_10360_out0;
assign v$STORE$PCOUNTER_2102_out0 = v$G6_11143_out0;
assign v$STORE$PCOUNTER_2103_out0 = v$G6_11144_out0;
assign v$_2146_out0 = { v$C1_10789_out0,v$_13253_out0 };
assign v$_2147_out0 = { v$C1_10790_out0,v$_13254_out0 };
assign v$MUX$ENABLE_2349_out0 = v$G16_3024_out0;
assign v$MULTI$INSTRUCTION_2451_out0 = v$MULTI$INSTRUCTION_13323_out0;
assign v$MULTI$INSTRUCTION_2452_out0 = v$MULTI$INSTRUCTION_13324_out0;
assign v$JMP_2668_out0 = v$JMP_7077_out0;
assign v$JMP_2669_out0 = v$JMP_7078_out0;
assign v$LOAD_3115_out0 = v$EQ2_7091_out0;
assign v$LOAD_3116_out0 = v$EQ2_7092_out0;
assign v$G26_4735_out0 = v$G23_2840_out0 && v$_2860_out0;
assign v$G26_4736_out0 = v$G23_2841_out0 && v$_2861_out0;
assign v$W$EN_6878_out0 = v$_10868_out1;
assign v$W$EN_6879_out0 = v$_10869_out1;
assign v$STALL_6910_out0 = v$STALL_427_out0;
assign v$STALL_6911_out0 = v$STALL_428_out0;
assign v$_7062_out0 = v$_10868_out0[6:0];
assign v$_7062_out1 = v$_10868_out0[7:1];
assign v$_7063_out0 = v$_10869_out0[6:0];
assign v$_7063_out1 = v$_10869_out0[7:1];
assign v$SUB$INSTRUCTION_7085_out0 = v$SUB$INSTRUCTION_11195_out0;
assign v$SUB$INSTRUCTION_7086_out0 = v$SUB$INSTRUCTION_11196_out0;
assign v$WEN1_7716_out0 = v$Wen1_10312_out0;
assign v$CMP_8646_out0 = v$CMP_3805_out0;
assign v$CMP_8647_out0 = v$CMP_3806_out0;
assign v$JMI_8679_out0 = v$JMI_88_out0;
assign v$JMI_8680_out0 = v$JMI_89_out0;
assign v$STP_10307_out0 = v$STP_10977_out0;
assign v$STP_10308_out0 = v$STP_10978_out0;
assign v$AD3_10482_out0 = v$MUX2_1145_out0;
assign v$AD3_10483_out0 = v$MUX2_1146_out0;
assign v$UART_10516_out0 = v$UART_10825_out0;
assign v$UART_10517_out0 = v$UART_10826_out0;
assign v$done$receiving_10604_out0 = v$BYTERECEIVED_11197_out0;
assign v$SR_10607_out0 = v$MUX1_534_out0;
assign v$SR_10608_out0 = v$MUX1_535_out0;
assign v$SBC_11051_out0 = v$SBC_4825_out0;
assign v$SBC_11052_out0 = v$SBC_4826_out0;
assign v$STP_11240_out0 = v$STP_10467_out0;
assign v$STP_11241_out0 = v$STP_10468_out0;
assign v$SUB_12247_out0 = v$SUB_2957_out0;
assign v$SUB_12248_out0 = v$SUB_2958_out0;
assign v$AD3_13272_out0 = v$MUX2_1145_out0;
assign v$AD3_13273_out0 = v$MUX2_1146_out0;
assign v$WEN0_13300_out0 = v$WEN0_2646_out0;
assign v$JEQ_13560_out0 = v$JEQ_4445_out0;
assign v$JEQ_13561_out0 = v$JEQ_4446_out0;
assign v$G1_13776_out0 = v$G2_2891_out0 || v$EXEC2_3241_out0;
assign v$G1_13777_out0 = v$G2_2892_out0 || v$EXEC2_3242_out0;
assign v$LOAD_231_out0 = v$LOAD_3115_out0;
assign v$LOAD_232_out0 = v$LOAD_3116_out0;
assign v$ROR_282_out0 = v$SR_542_out0 == 2'h3;
assign v$ROR_283_out0 = v$SR_543_out0 == 2'h3;
assign v$G6_327_out0 = v$C_3197_out0 && v$ADC_1821_out0;
assign v$G6_328_out0 = v$C_3198_out0 && v$ADC_1822_out0;
assign v$G9_407_out0 = ! v$W$EN_6878_out0;
assign v$G9_408_out0 = ! v$W$EN_6879_out0;
assign v$G9_411_out0 = ((v$AND_13556_out0 && !v$TST_409_out0) || (!v$AND_13556_out0) && v$TST_409_out0);
assign v$G9_412_out0 = ((v$AND_13557_out0 && !v$TST_410_out0) || (!v$AND_13557_out0) && v$TST_410_out0);
assign v$LSR_418_out0 = v$SR_371_out0 == 2'h1;
assign v$LSR_419_out0 = v$SR_372_out0 == 2'h1;
assign v$G5_454_out0 = v$STORE_1195_out0 && v$EXEC1_20_out0;
assign v$G5_455_out0 = v$STORE_1196_out0 && v$EXEC1_21_out0;
assign v$RD_501_out0 = v$DOUT1_1207_out0;
assign v$RD_502_out0 = v$DOUT1_1208_out0;
assign v$STORE_540_out0 = v$STORE_1195_out0;
assign v$STORE_541_out0 = v$STORE_1196_out0;
assign v$ROR_544_out0 = v$SR_371_out0 == 2'h3;
assign v$ROR_545_out0 = v$SR_372_out0 == 2'h3;
assign v$LSR_1174_out0 = v$SR_542_out0 == 2'h1;
assign v$LSR_1175_out0 = v$SR_543_out0 == 2'h1;
assign v$G9_1671_out0 = ! v$STALL_6910_out0;
assign v$G9_1672_out0 = ! v$STALL_6911_out0;
assign v$LSL_1861_out0 = v$SR_542_out0 == 2'h0;
assign v$LSL_1862_out0 = v$SR_543_out0 == 2'h0;
assign v$G2_1887_out0 = v$W$EN_6878_out0 && v$EXEC1_20_out0;
assign v$G2_1888_out0 = v$W$EN_6879_out0 && v$EXEC1_21_out0;
assign v$MUX1_2409_out0 = v$C_379_out0 ? v$_2146_out0 : v$BIN_5853_out0;
assign v$MUX1_2410_out0 = v$C_380_out0 ? v$_2147_out0 : v$BIN_5854_out0;
assign v$LSL_2842_out0 = v$SR_10607_out0 == 2'h0;
assign v$LSL_2843_out0 = v$SR_10608_out0 == 2'h0;
assign v$STORE$pccounter_2883_out0 = v$STORE$PCOUNTER_2102_out0;
assign v$STORE$pccounter_2884_out0 = v$STORE$PCOUNTER_2103_out0;
assign v$G3_2903_out0 = v$LOAD_3115_out0 && v$EXEC2_7181_out0;
assign v$G3_2904_out0 = v$LOAD_3116_out0 && v$EXEC2_7182_out0;
assign v$G1_3018_out0 = v$SBC_11051_out0 && v$C_3197_out0;
assign v$G1_3019_out0 = v$SBC_11052_out0 && v$C_3198_out0;
assign v$LSL_3047_out0 = v$SR_371_out0 == 2'h0;
assign v$LSL_3048_out0 = v$SR_372_out0 == 2'h0;
assign v$LSL_3182_out0 = v$SR_1956_out0 == 2'h0;
assign v$LSL_3183_out0 = v$SR_1957_out0 == 2'h0;
assign v$ROR_3286_out0 = v$SR_10607_out0 == 2'h3;
assign v$ROR_3287_out0 = v$SR_10608_out0 == 2'h3;
assign v$ROR_3288_out0 = v$SR_1956_out0 == 2'h3;
assign v$ROR_3289_out0 = v$SR_1957_out0 == 2'h3;
assign v$UART_3893_out0 = v$UART_10516_out0;
assign v$UART_3894_out0 = v$UART_10517_out0;
assign v$G5_4477_out0 = v$SUB_12247_out0 || v$CMP_8646_out0;
assign v$G5_4478_out0 = v$SUB_12248_out0 || v$CMP_8647_out0;
assign v$G4_4738_out0 = ((v$SBC_11051_out0 && !v$ADC_1821_out0) || (!v$SBC_11051_out0) && v$ADC_1821_out0);
assign v$G4_4739_out0 = ((v$SBC_11052_out0 && !v$ADC_1822_out0) || (!v$SBC_11052_out0) && v$ADC_1822_out0);
assign v$G29_5834_out0 = v$G26_4735_out0 || v$G27_9793_out0;
assign v$G29_5835_out0 = v$G26_4736_out0 || v$G27_9794_out0;
assign v$LSR_6912_out0 = v$SR_1956_out0 == 2'h1;
assign v$LSR_6913_out0 = v$SR_1957_out0 == 2'h1;
assign v$G3_8665_out0 = ((v$SUB_12247_out0 && !v$CMP_8646_out0) || (!v$SUB_12247_out0) && v$CMP_8646_out0);
assign v$G3_8666_out0 = ((v$SUB_12248_out0 && !v$CMP_8647_out0) || (!v$SUB_12248_out0) && v$CMP_8647_out0);
assign v$AD3_8671_out0 = v$AD3_13272_out0;
assign v$AD3_8672_out0 = v$AD3_13273_out0;
assign v$ASR_8754_out0 = v$SR_1956_out0 == 2'h2;
assign v$ASR_8755_out0 = v$SR_1957_out0 == 2'h2;
assign v$G18_8799_out0 = !(v$ENABLE_2018_out0 || v$Q7_6888_out0);
assign v$STALL_10281_out0 = v$STALL_1758_out0;
assign v$STALL_10282_out0 = v$STALL_1759_out0;
assign v$G4_10283_out0 = v$G5_10914_out0 && v$STALL_6910_out0;
assign v$G4_10284_out0 = v$G5_10915_out0 && v$STALL_6911_out0;
assign v$G19_10327_out0 = ! v$STP_11240_out0;
assign v$G19_10328_out0 = ! v$STP_11241_out0;
assign v$ASR_10366_out0 = v$SR_542_out0 == 2'h2;
assign v$ASR_10367_out0 = v$SR_543_out0 == 2'h2;
assign v$RX$DONE$RECEIVING_10484_out0 = v$done$receiving_10604_out0;
assign v$_10490_out0 = v$_7062_out0[5:0];
assign v$_10490_out1 = v$_7062_out0[6:1];
assign v$_10491_out0 = v$_7063_out0[5:0];
assign v$_10491_out1 = v$_7063_out0[6:1];
assign v$ASR_10566_out0 = v$SR_371_out0 == 2'h2;
assign v$ASR_10567_out0 = v$SR_372_out0 == 2'h2;
assign v$P_10682_out0 = v$_7062_out1;
assign v$P_10683_out0 = v$_7063_out1;
assign v$G17_10710_out0 = v$MUX$ENABLE_2349_out0 && v$G18_567_out0;
assign v$WENMULTI_11206_out0 = v$G1_13776_out0;
assign v$WENMULTI_11207_out0 = v$G1_13777_out0;
assign v$G4_12243_out0 = v$G5_10441_out0 && v$G3_17_out0;
assign v$G4_12244_out0 = v$G5_10442_out0 && v$G3_18_out0;
assign v$MULTI$INSTRUCTION_13308_out0 = v$MULTI$INSTRUCTION_619_out0;
assign v$MULTI$INSTRUCTION_13309_out0 = v$MULTI$INSTRUCTION_620_out0;
assign v$LSR_13331_out0 = v$SR_10607_out0 == 2'h1;
assign v$LSR_13332_out0 = v$SR_10608_out0 == 2'h1;
assign v$G11_13439_out0 = v$G20_598_out0 || v$STP_11240_out0;
assign v$G11_13440_out0 = v$G20_599_out0 || v$STP_11241_out0;
assign v$RM_13597_out0 = v$DOUT2_1733_out0;
assign v$RM_13598_out0 = v$DOUT2_1734_out0;
assign v$ASR_13713_out0 = v$SR_10607_out0 == 2'h2;
assign v$ASR_13714_out0 = v$SR_10608_out0 == 2'h2;
assign v$RM_13750_out0 = v$DOUT2_1733_out0;
assign v$RM_13751_out0 = v$DOUT2_1734_out0;
assign v$G30_184_out0 = v$G2_1888_out0 && v$STALL$DUAL$CORE_12235_out0;
assign v$_1140_out0 = v$_10490_out0[1:0];
assign v$_1140_out1 = v$_10490_out0[5:4];
assign v$_1141_out0 = v$_10491_out0[1:0];
assign v$_1141_out1 = v$_10491_out0[5:4];
assign v$G1_1191_out0 = ! v$_10490_out1;
assign v$G1_1192_out0 = ! v$_10491_out1;
assign v$G8_1765_out0 = v$G7_1684_out0 || v$G4_10283_out0;
assign v$G8_1766_out0 = v$G7_1685_out0 || v$G4_10284_out0;
assign v$G22_1900_out0 = v$G11_13440_out0 && v$STALL$DUAL$CORE_4696_out0;
assign v$WEN$MULTI_2388_out0 = v$WENMULTI_11206_out0;
assign v$WEN$MULTI_2389_out0 = v$WENMULTI_11207_out0;
assign v$G11_2626_out0 = v$G5_10914_out0 && v$G9_1671_out0;
assign v$G11_2627_out0 = v$G5_10915_out0 && v$G9_1672_out0;
assign v$RDOUT_2787_out0 = v$RD_501_out0;
assign v$RDOUT_2788_out0 = v$RD_502_out0;
assign v$LOAD_2899_out0 = v$LOAD_231_out0;
assign v$LOAD_2900_out0 = v$LOAD_232_out0;
assign v$DONE$RECEIVING_3084_out0 = v$RX$DONE$RECEIVING_10484_out0;
assign v$RXBYTERECEIVED_3269_out0 = v$RX$DONE$RECEIVING_10484_out0;
assign v$G21_3808_out0 = v$G18_8799_out0 || v$G22_10983_out0;
assign v$RD_3891_out0 = v$RD_501_out0;
assign v$RD_3892_out0 = v$RD_502_out0;
assign v$OP1_3899_out0 = v$RD_501_out0;
assign v$OP1_3900_out0 = v$RD_502_out0;
assign v$G8_4453_out0 = v$G1_3018_out0 || v$G6_327_out0;
assign v$G8_4454_out0 = v$G1_3019_out0 || v$G6_328_out0;
assign v$G7_4474_out0 = v$P_10682_out0 && v$EXEC1_20_out0;
assign v$G7_4475_out0 = v$P_10683_out0 && v$EXEC1_21_out0;
assign v$G10_4479_out0 = v$EXEC2_7181_out0 && v$P_10682_out0;
assign v$G10_4480_out0 = v$EXEC2_7182_out0 && v$P_10683_out0;
assign v$RM_4537_out0 = v$RM_13750_out0;
assign v$RM_4538_out0 = v$RM_13751_out0;
assign v$STORE$WEN_4544_out0 = v$STORE$pccounter_2883_out0;
assign v$STORE$WEN_4545_out0 = v$STORE$pccounter_2884_out0;
assign v$EN_4593_out0 = v$G29_5834_out0;
assign v$EN_4594_out0 = v$G29_5835_out0;
assign v$G24_4780_out0 = ! v$G17_10710_out0;
assign v$G5_7106_out0 = v$MULTI$INSTRUCTION_13308_out0 || v$DIV$INSTRUCTION_4614_out0;
assign v$G5_7107_out0 = v$MULTI$INSTRUCTION_13309_out0 || v$DIV$INSTRUCTION_4615_out0;
assign v$RM_8731_out0 = v$RM_13750_out0;
assign v$RM_8732_out0 = v$RM_13751_out0;
assign v$MUX1_8813_out0 = v$C_8653_out0 ? v$KEXTEND_13329_out0 : v$RM_13597_out0;
assign v$MUX1_8814_out0 = v$C_8654_out0 ? v$KEXTEND_13330_out0 : v$RM_13598_out0;
assign v$MUX10_10395_out0 = v$MULTI$INSTRUCTION_13308_out0 ? v$C13_405_out0 : v$C12_2113_out0;
assign v$MUX10_10396_out0 = v$MULTI$INSTRUCTION_13309_out0 ? v$C13_406_out0 : v$C12_2114_out0;
assign v$RAMWEN_10701_out0 = v$G5_454_out0;
assign v$RAMWEN_10702_out0 = v$G5_455_out0;
assign v$B_10793_out0 = v$MUX1_2409_out0;
assign v$B_10794_out0 = v$MUX1_2410_out0;
assign v$STORE_10831_out0 = v$STORE_540_out0;
assign v$STORE_10832_out0 = v$STORE_541_out0;
assign v$WENALU_10866_out0 = v$G4_12243_out0;
assign v$WENALU_10867_out0 = v$G4_12244_out0;
assign v$UART_11128_out0 = v$UART_3893_out0;
assign v$UART_11129_out0 = v$UART_3894_out0;
assign v$G2_11134_out0 = ((v$ADD_11193_out0 && !v$G3_8665_out0) || (!v$ADD_11193_out0) && v$G3_8665_out0);
assign v$G2_11135_out0 = ((v$ADD_11194_out0 && !v$G3_8666_out0) || (!v$ADD_11194_out0) && v$G3_8666_out0);
assign v$G11_11165_out0 = v$G5_4477_out0 || v$SBC_11051_out0;
assign v$G11_11166_out0 = v$G5_4478_out0 || v$SBC_11052_out0;
assign v$RM_11167_out0 = v$RM_13750_out0;
assign v$RM_11168_out0 = v$RM_13751_out0;
assign v$G4_13702_out0 = ! v$MULTI$INSTRUCTION_13308_out0;
assign v$G4_13703_out0 = ! v$MULTI$INSTRUCTION_13309_out0;
assign v$EN$STALL_13747_out0 = v$G17_10710_out0;
assign v$RXBYTERECEIVED_91_out0 = v$RXBYTERECEIVED_3269_out0;
assign v$SEL6_103_out0 = v$RM_11167_out0[9:0];
assign v$SEL6_104_out0 = v$RM_11168_out0[9:0];
assign v$G10_130_out0 = v$G8_4453_out0 || v$G5_4477_out0;
assign v$G10_131_out0 = v$G8_4454_out0 || v$G5_4478_out0;
assign v$G7_169_out0 = ((v$G2_11134_out0 && !v$G4_4738_out0) || (!v$G2_11134_out0) && v$G4_4738_out0);
assign v$G7_170_out0 = ((v$G2_11135_out0 && !v$G4_4739_out0) || (!v$G2_11135_out0) && v$G4_4739_out0);
assign v$_186_out0 = v$B_10793_out0[3:3];
assign v$_187_out0 = v$B_10794_out0[3:3];
assign v$G4_220_out0 = v$G30_184_out0 || v$G3_2904_out0;
assign v$_413_out0 = v$B_10793_out0[1:1];
assign v$_414_out0 = v$B_10794_out0[1:1];
assign v$_1728_out0 = v$B_10793_out0[0:0];
assign v$_1729_out0 = v$B_10794_out0[0:0];
assign v$WENRAM_2326_out0 = v$RAMWEN_10701_out0;
assign v$WENRAM_2327_out0 = v$RAMWEN_10702_out0;
assign v$G18_2407_out0 = v$G16_2310_out0 && v$G8_1765_out0;
assign v$G18_2408_out0 = v$G16_2311_out0 && v$G8_1766_out0;
assign v$RM_2432_out0 = v$RM_8731_out0;
assign v$RM_2433_out0 = v$RM_8732_out0;
assign v$SEL3_2615_out0 = v$RD_3891_out0[15:15];
assign v$SEL3_2616_out0 = v$RD_3892_out0[15:15];
assign v$G8_2623_out0 = v$G9_407_out0 && v$G10_4479_out0;
assign v$G8_2624_out0 = v$G9_408_out0 && v$G10_4480_out0;
assign v$SUB_2910_out0 = v$G22_1900_out0;
assign v$SEL1_2917_out0 = v$RD_3891_out0[14:10];
assign v$SEL1_2918_out0 = v$RD_3892_out0[14:10];
assign v$OP1_2979_out0 = v$OP1_3899_out0;
assign v$OP1_2980_out0 = v$OP1_3900_out0;
assign v$G23_3083_out0 = v$WEN1_7716_out0 && v$G24_4780_out0;
assign v$SUB_4616_out0 = v$G11_11165_out0;
assign v$SUB_4618_out0 = v$G11_11166_out0;
assign v$M_4701_out0 = v$_1140_out0;
assign v$M_4702_out0 = v$_1141_out0;
assign v$DONE$RECEIVING_5857_out0 = v$DONE$RECEIVING_3084_out0;
assign v$LOAD_7110_out0 = v$LOAD_2899_out0;
assign v$LOAD_7111_out0 = v$LOAD_2900_out0;
assign v$SEL4_7636_out0 = v$RM_11167_out0[15:15];
assign v$SEL4_7637_out0 = v$RM_11168_out0[15:15];
assign v$N_7642_out0 = v$_1140_out1;
assign v$N_7643_out0 = v$_1141_out1;
assign v$WENALU_8659_out0 = v$WENALU_10866_out0;
assign v$WENALU_8660_out0 = v$WENALU_10867_out0;
assign v$SEL5_8767_out0 = v$RD_3891_out0[9:0];
assign v$SEL5_8768_out0 = v$RD_3892_out0[9:0];
assign v$REGISTER$OUT_10268_out0 = v$RDOUT_2787_out0;
assign v$REGISTER$OUT_10269_out0 = v$RDOUT_2788_out0;
assign v$G12_10321_out0 = v$G11_2626_out0 && v$G2_6791_out0;
assign v$G12_10322_out0 = v$G11_2627_out0 && v$G2_6792_out0;
assign v$EN$STALL_10344_out0 = v$EN$STALL_13747_out0;
assign v$WEN$MULTI_10381_out0 = v$WEN$MULTI_2388_out0;
assign v$WEN$MULTI_10382_out0 = v$WEN$MULTI_2389_out0;
assign v$U_10469_out0 = v$G1_1191_out0;
assign v$U_10470_out0 = v$G1_1192_out0;
assign v$_10785_out0 = v$B_10793_out0[2:2];
assign v$_10786_out0 = v$B_10794_out0[2:2];
assign v$IN_11258_out0 = v$MUX1_8813_out0;
assign v$IN_11259_out0 = v$MUX1_8814_out0;
assign v$STORE_13298_out0 = v$STORE_10831_out0;
assign v$STORE_13299_out0 = v$STORE_10832_out0;
assign v$SEL2_13327_out0 = v$RM_11167_out0[14:10];
assign v$SEL2_13328_out0 = v$RM_11168_out0[14:10];
assign v$RM_13508_out0 = v$RM_4537_out0;
assign v$RM_13509_out0 = v$RM_4538_out0;
assign v$WEN$MULTI_35_out0 = v$WEN$MULTI_10381_out0;
assign v$WEN$MULTI_36_out0 = v$WEN$MULTI_10382_out0;
assign v$IN_98_out0 = v$IN_11258_out0;
assign v$IN_99_out0 = v$IN_11259_out0;
assign v$STORE_221_out0 = v$STORE_13298_out0;
assign v$STORE_222_out0 = v$STORE_13299_out0;
assign v$G5_230_out0 = ((v$_3271_out0 && !v$SUB_2910_out0) || (!v$_3271_out0) && v$SUB_2910_out0);
assign v$RAM$IN_233_out0 = v$REGISTER$OUT_10268_out0;
assign v$RAM$IN_234_out0 = v$REGISTER$OUT_10269_out0;
assign v$RD$SIGN_285_out0 = v$SEL3_2615_out0;
assign v$RD$SIGN_286_out0 = v$SEL3_2616_out0;
assign v$G10_1755_out0 = v$G6_2905_out0 || v$G12_10321_out0;
assign v$G10_1756_out0 = v$G6_2906_out0 || v$G12_10322_out0;
assign v$RD$SIG_1769_out0 = v$SEL5_8767_out0;
assign v$RD$SIG_1770_out0 = v$SEL5_8768_out0;
assign v$G17_1903_out0 = v$RXBYTERECEIVED_91_out0 && v$Q1_3993_out0;
assign v$G8_2025_out0 = ((v$_172_out0 && !v$SUB_2910_out0) || (!v$_172_out0) && v$SUB_2910_out0);
assign v$OP1_2060_out0 = v$OP1_2979_out0;
assign v$OP1_2061_out0 = v$OP1_2980_out0;
assign v$EN_2330_out0 = v$_1728_out0;
assign v$EN_2331_out0 = v$_1729_out0;
assign v$G9_2333_out0 = ((v$_2269_out0 && !v$SUB_2910_out0) || (!v$_2269_out0) && v$SUB_2910_out0);
assign v$G6_2417_out0 = ((v$_2023_out0 && !v$SUB_2910_out0) || (!v$_2023_out0) && v$SUB_2910_out0);
assign v$EN_2445_out0 = v$_186_out0;
assign v$EN_2446_out0 = v$_187_out0;
assign v$OP2$EXP_2548_out0 = v$SEL2_13327_out0;
assign v$OP2$EXP_2549_out0 = v$SEL2_13328_out0;
assign v$G11_2551_out0 = ((v$_61_out0 && !v$SUB_2910_out0) || (!v$_61_out0) && v$SUB_2910_out0);
assign v$G3_2622_out0 = ((v$_288_out0 && !v$SUB_2910_out0) || (!v$_288_out0) && v$SUB_2910_out0);
assign v$G10_2633_out0 = ((v$_11243_out0 && !v$SUB_2910_out0) || (!v$_11243_out0) && v$SUB_2910_out0);
assign v$_3035_out0 = v$RM_13508_out0[11:0];
assign v$_3035_out1 = v$RM_13508_out0[15:4];
assign v$_3036_out0 = v$RM_13509_out0[11:0];
assign v$_3036_out1 = v$RM_13509_out0[15:4];
assign v$G2_3240_out0 = ((v$_3124_out0 && !v$SUB_2910_out0) || (!v$_3124_out0) && v$SUB_2910_out0);
assign v$G19_3860_out0 = v$RXBYTERECEIVED_91_out0 || v$Q1_3993_out0;
assign v$SUB_4617_out0 = v$U_10469_out0;
assign v$SUB_4619_out0 = v$U_10470_out0;
assign v$WENRAM_4650_out0 = v$WENRAM_2326_out0;
assign v$WENRAM_4651_out0 = v$WENRAM_2327_out0;
assign v$G12_4700_out0 = ((v$_1876_out0 && !v$SUB_2910_out0) || (!v$_1876_out0) && v$SUB_2910_out0);
assign v$G7_4822_out0 = ((v$_13397_out0 && !v$SUB_2910_out0) || (!v$_13397_out0) && v$SUB_2910_out0);
assign v$byte$ready_5843_out0 = v$DONE$RECEIVING_5857_out0;
assign v$LOAD_8765_out0 = v$LOAD_7110_out0;
assign v$LOAD_8766_out0 = v$LOAD_7111_out0;
assign v$RD$EXP_8846_out0 = v$SEL1_2917_out0;
assign v$RD$EXP_8847_out0 = v$SEL1_2918_out0;
assign v$EN_10474_out0 = v$_413_out0;
assign v$EN_10475_out0 = v$_414_out0;
assign v$G1_10478_out0 = ((v$_13563_out0 && !v$SUB_2910_out0) || (!v$_13563_out0) && v$SUB_2910_out0);
assign v$G21_10788_out0 = v$G23_3083_out0 || v$WEN0_13300_out0;
assign v$OP2$SIGN_10839_out0 = v$SEL4_7636_out0;
assign v$OP2$SIGN_10840_out0 = v$SEL4_7637_out0;
assign v$_11229_out0 = { v$N_7642_out0,v$C1_3210_out0 };
assign v$_11230_out0 = { v$N_7643_out0,v$C1_3211_out0 };
assign v$G4_12239_out0 = ((v$_180_out0 && !v$SUB_2910_out0) || (!v$_180_out0) && v$SUB_2910_out0);
assign v$EN_13181_out0 = v$_10785_out0;
assign v$EN_13182_out0 = v$_10786_out0;
assign v$G6_13258_out0 = v$G8_2623_out0 || v$G7_4474_out0;
assign v$G6_13259_out0 = v$G8_2624_out0 || v$G7_4475_out0;
assign v$OP2$SIG_13301_out0 = v$SEL6_103_out0;
assign v$OP2$SIG_13302_out0 = v$SEL6_104_out0;
assign v$STALL$DUAL$CORE_13617_out0 = v$EN$STALL_10344_out0;
assign v$WENLDST_13756_out0 = v$G4_220_out0;
assign v$OP2$EXP_536_out0 = v$OP2$EXP_2548_out0;
assign v$OP2$EXP_537_out0 = v$OP2$EXP_2549_out0;
assign v$_1708_out0 = { v$G1_10478_out0,v$G2_3240_out0 };
assign v$SIG$RM_1767_out0 = v$OP2$SIG_13301_out0;
assign v$SIG$RM_1768_out0 = v$OP2$SIG_13302_out0;
assign v$RD$SIGN_2405_out0 = v$RD$SIGN_285_out0;
assign v$RD$SIGN_2406_out0 = v$RD$SIGN_286_out0;
assign v$WENLDST_2683_out0 = v$WENLDST_13756_out0;
assign v$WEN_3204_out0 = v$G21_10788_out0;
assign v$LOAD_3949_out0 = v$LOAD_8765_out0;
assign v$LOAD_3950_out0 = v$LOAD_8766_out0;
assign v$RD$EXP_3951_out0 = v$RD$EXP_8846_out0;
assign v$RD$EXP_3952_out0 = v$RD$EXP_8847_out0;
assign v$G2_4467_out0 = ! v$STALL$DUAL$CORE_13617_out0;
assign v$EXP$RM_4743_out0 = v$OP2$EXP_2548_out0;
assign v$EXP$RM_4744_out0 = v$OP2$EXP_2549_out0;
assign v$_4831_out0 = v$IN_98_out0[14:0];
assign v$_4831_out1 = v$IN_98_out0[15:1];
assign v$_4832_out0 = v$IN_99_out0[14:0];
assign v$_4832_out1 = v$IN_99_out0[15:1];
assign v$EXP$RD_5855_out0 = v$RD$EXP_8846_out0;
assign v$EXP$RD_5856_out0 = v$RD$EXP_8847_out0;
assign v$A_10275_out0 = v$OP1_2060_out0;
assign v$A_10277_out0 = v$OP1_2061_out0;
assign v$BYTE$READY_11173_out0 = v$byte$ready_5843_out0;
assign v$OP2$SIGN_11208_out0 = v$OP2$SIGN_10839_out0;
assign v$OP2$SIGN_11209_out0 = v$OP2$SIGN_10840_out0;
assign v$A_11251_out0 = v$_11229_out0;
assign v$A_11253_out0 = v$_11230_out0;
assign v$SIG$RD_11298_out0 = v$RD$SIG_1769_out0;
assign v$SIG$RD_11299_out0 = v$RD$SIG_1770_out0;
assign v$G14_13268_out0 = v$G10_1755_out0 || v$G13_7083_out0;
assign v$G14_13269_out0 = v$G10_1756_out0 || v$G13_7084_out0;
assign v$UNUSED_13431_out0 = v$_3035_out1;
assign v$UNUSED_13432_out0 = v$_3036_out1;
assign v$IN_13788_out0 = v$IN_98_out0;
assign v$IN_13789_out0 = v$IN_99_out0;
assign v$_1_out0 = v$A_10275_out0[4:4];
assign v$_3_out0 = v$A_10277_out0[4:4];
assign v$_78_out0 = v$A_11251_out0[3:3];
assign v$_80_out0 = v$A_11253_out0[3:3];
assign v$_193_out0 = v$A_11251_out0[15:15];
assign v$_195_out0 = v$A_11253_out0[15:15];
assign v$G1_289_out0 = ((v$OP2$SIGN_11208_out0 && !v$SUB$INSTRUCTION_7085_out0) || (!v$OP2$SIGN_11208_out0) && v$SUB$INSTRUCTION_7085_out0);
assign v$G1_290_out0 = ((v$OP2$SIGN_11209_out0 && !v$SUB$INSTRUCTION_7086_out0) || (!v$OP2$SIGN_11209_out0) && v$SUB$INSTRUCTION_7086_out0);
assign v$_322_out0 = v$A_11251_out0[0:0];
assign v$_324_out0 = v$A_11253_out0[0:0];
assign v$_330_out0 = v$A_11251_out0[9:9];
assign v$_332_out0 = v$A_11253_out0[9:9];
assign v$WENLS_601_out0 = v$WENLDST_2683_out0;
assign v$_1693_out0 = v$A_10275_out0[5:5];
assign v$_1695_out0 = v$A_10277_out0[5:5];
assign v$_1748_out0 = v$A_10275_out0[11:11];
assign v$_1750_out0 = v$A_10277_out0[11:11];
assign v$_1894_out0 = v$A_10275_out0[0:0];
assign v$_1896_out0 = v$A_10277_out0[0:0];
assign v$_2094_out0 = v$A_11251_out0[13:13];
assign v$_2096_out0 = v$A_11253_out0[13:13];
assign v$_2151_out0 = v$A_10275_out0[2:2];
assign v$_2153_out0 = v$A_10277_out0[2:2];
assign v$WEN_2154_out0 = v$WEN_3204_out0;
assign v$_2387_out0 = { v$_1708_out0,v$G3_2622_out0 };
assign v$_2419_out0 = v$A_11251_out0[6:6];
assign v$_2421_out0 = v$A_11253_out0[6:6];
assign v$RD$EXP_2601_out0 = v$RD$EXP_3951_out0;
assign v$RD$EXP_2602_out0 = v$RD$EXP_3952_out0;
assign v$_2761_out0 = v$A_10275_out0[15:15];
assign v$_2763_out0 = v$A_10277_out0[15:15];
assign v$_2876_out0 = v$A_10275_out0[12:12];
assign v$_2878_out0 = v$A_10277_out0[12:12];
assign v$_2880_out0 = v$A_10275_out0[3:3];
assign v$_2882_out0 = v$A_10277_out0[3:3];
assign v$_3120_out0 = v$A_11251_out0[14:14];
assign v$_3122_out0 = v$A_11253_out0[14:14];
assign v$STALL$DUAL$CORE_3127_out0 = v$G2_4467_out0;
assign v$_3248_out0 = v$A_10275_out0[8:8];
assign v$_3250_out0 = v$A_10277_out0[8:8];
assign v$_3283_out0 = v$A_11251_out0[2:2];
assign v$_3285_out0 = v$A_11253_out0[2:2];
assign v$_4598_out0 = v$A_10275_out0[10:10];
assign v$_4600_out0 = v$A_10277_out0[10:10];
assign v$_4712_out0 = v$A_10275_out0[13:13];
assign v$_4714_out0 = v$A_10277_out0[13:13];
assign v$BYTE$READY_7022_out0 = v$BYTE$READY_11173_out0;
assign v$_7179_out0 = { v$C1_604_out0,v$_4831_out0 };
assign v$_7180_out0 = { v$C1_605_out0,v$_4832_out0 };
assign v$_8749_out0 = v$A_11251_out0[8:8];
assign v$_8751_out0 = v$A_11253_out0[8:8];
assign v$MUX3_8818_out0 = v$IR15_2465_out0 ? v$WENALU_8660_out0 : v$WENLDST_2683_out0;
assign v$_8828_out0 = v$A_11251_out0[7:7];
assign v$_8830_out0 = v$A_11253_out0[7:7];
assign v$_8849_out0 = v$A_10275_out0[14:14];
assign v$_8851_out0 = v$A_10277_out0[14:14];
assign v$EQ2_10347_out0 = v$EXP$RM_4743_out0 == 5'h0;
assign v$EQ2_10348_out0 = v$EXP$RM_4744_out0 == 5'h0;
assign v$_10378_out0 = v$A_11251_out0[5:5];
assign v$_10380_out0 = v$A_11253_out0[5:5];
assign v$OP2$EXP_10383_out0 = v$OP2$EXP_536_out0;
assign v$OP2$EXP_10384_out0 = v$OP2$EXP_537_out0;
assign v$_10386_out0 = v$A_11251_out0[1:1];
assign v$_10388_out0 = v$A_11253_out0[1:1];
assign v$_10696_out0 = v$A_11251_out0[4:4];
assign v$_10698_out0 = v$A_11253_out0[4:4];
assign v$_10778_out0 = v$A_11251_out0[12:12];
assign v$_10780_out0 = v$A_11253_out0[12:12];
assign v$_10863_out0 = v$A_11251_out0[10:10];
assign v$_10865_out0 = v$A_11253_out0[10:10];
assign v$_11057_out0 = { v$G14_13268_out0,v$G18_2407_out0 };
assign v$_11058_out0 = { v$G14_13269_out0,v$G18_2408_out0 };
assign v$_11150_out0 = v$A_10275_out0[6:6];
assign v$_11152_out0 = v$A_10277_out0[6:6];
assign v$UNNOTUSED_11220_out0 = v$_4831_out1;
assign v$UNNOTUSED_11221_out0 = v$_4832_out1;
assign v$_13385_out0 = v$A_10275_out0[7:7];
assign v$_13387_out0 = v$A_10277_out0[7:7];
assign v$EQ1_13433_out0 = v$EXP$RD_5855_out0 == 5'h0;
assign v$EQ1_13434_out0 = v$EXP$RD_5856_out0 == 5'h0;
assign v$_13513_out0 = v$A_10275_out0[1:1];
assign v$_13515_out0 = v$A_10277_out0[1:1];
assign v$_13553_out0 = v$A_11251_out0[11:11];
assign v$_13555_out0 = v$A_11253_out0[11:11];
assign v$_13628_out0 = v$A_10275_out0[9:9];
assign v$_13630_out0 = v$A_10277_out0[9:9];
assign v$MUX1_31_out0 = v$LSL_3182_out0 ? v$_7179_out0 : v$IN_13788_out0;
assign v$MUX1_32_out0 = v$LSL_3183_out0 ? v$_7180_out0 : v$IN_13789_out0;
assign v$G3_207_out0 = ((v$_3283_out0 && !v$SUB_4617_out0) || (!v$_3283_out0) && v$SUB_4617_out0);
assign v$G3_209_out0 = ((v$_3285_out0 && !v$SUB_4619_out0) || (!v$_3285_out0) && v$SUB_4619_out0);
assign v$D_623_out0 = v$_11057_out0;
assign v$D_624_out0 = v$_11058_out0;
assign v$G1_646_out0 = ! v$EQ1_13433_out0;
assign v$G1_647_out0 = ! v$EQ1_13434_out0;
assign v$G8_1216_out0 = ((v$_8828_out0 && !v$SUB_4617_out0) || (!v$_8828_out0) && v$SUB_4617_out0);
assign v$G8_1218_out0 = ((v$_8830_out0 && !v$SUB_4619_out0) || (!v$_8830_out0) && v$SUB_4619_out0);
assign v$STALL$DUAL$CORE_1738_out0 = v$STALL$DUAL$CORE_3127_out0;
assign v$EQ2_1753_out0 = v$OP2$EXP_10383_out0 == 5'h0;
assign v$EQ2_1754_out0 = v$OP2$EXP_10384_out0 == 5'h0;
assign v$G15_1815_out0 = ((v$_3120_out0 && !v$SUB_4617_out0) || (!v$_3120_out0) && v$SUB_4617_out0);
assign v$G15_1817_out0 = ((v$_3122_out0 && !v$SUB_4619_out0) || (!v$_3122_out0) && v$SUB_4619_out0);
assign v$EQ1_2597_out0 = v$RD$EXP_2601_out0 == 5'h0;
assign v$EQ1_2598_out0 = v$RD$EXP_2602_out0 == 5'h0;
assign v$G7_2780_out0 = ((v$_2419_out0 && !v$SUB_4617_out0) || (!v$_2419_out0) && v$SUB_4617_out0);
assign v$G7_2782_out0 = ((v$_2421_out0 && !v$SUB_4619_out0) || (!v$_2421_out0) && v$SUB_4619_out0);
assign v$_2969_out0 = { v$_2387_out0,v$G4_12239_out0 };
assign v$STALL$DUAL$CORE_3264_out0 = v$STALL$DUAL$CORE_3127_out0;
assign v$G12_3346_out0 = ((v$_13553_out0 && !v$SUB_4617_out0) || (!v$_13553_out0) && v$SUB_4617_out0);
assign v$G12_3348_out0 = ((v$_13555_out0 && !v$SUB_4619_out0) || (!v$_13555_out0) && v$SUB_4619_out0);
assign v$G14_4534_out0 = ((v$_2094_out0 && !v$SUB_4617_out0) || (!v$_2094_out0) && v$SUB_4617_out0);
assign v$G14_4536_out0 = ((v$_2096_out0 && !v$SUB_4619_out0) || (!v$_2096_out0) && v$SUB_4619_out0);
assign v$G13_4706_out0 = ((v$_10778_out0 && !v$SUB_4617_out0) || (!v$_10778_out0) && v$SUB_4617_out0);
assign v$G13_4708_out0 = ((v$_10780_out0 && !v$SUB_4619_out0) || (!v$_10780_out0) && v$SUB_4619_out0);
assign v$G2_7015_out0 = ! v$EQ2_10347_out0;
assign v$G2_7016_out0 = ! v$EQ2_10348_out0;
assign v$G2_7026_out0 = ((v$_10386_out0 && !v$SUB_4617_out0) || (!v$_10386_out0) && v$SUB_4617_out0);
assign v$G2_7028_out0 = ((v$_10388_out0 && !v$SUB_4619_out0) || (!v$_10388_out0) && v$SUB_4619_out0);
assign v$MUX6_8758_out0 = v$MULTI$OPCODE_3021_out0 ? v$WEN$MULTI_2389_out0 : v$MUX3_8818_out0;
assign v$BYTE$READY_10559_out0 = v$BYTE$READY_7022_out0;
assign v$G5_10569_out0 = ((v$_10696_out0 && !v$SUB_4617_out0) || (!v$_10696_out0) && v$SUB_4617_out0);
assign v$G5_10571_out0 = ((v$_10698_out0 && !v$SUB_4619_out0) || (!v$_10698_out0) && v$SUB_4619_out0);
assign v$G4_10998_out0 = ((v$_78_out0 && !v$SUB_4617_out0) || (!v$_78_out0) && v$SUB_4617_out0);
assign v$G4_11000_out0 = ((v$_80_out0 && !v$SUB_4619_out0) || (!v$_80_out0) && v$SUB_4619_out0);
assign v$G16_11035_out0 = ((v$_193_out0 && !v$SUB_4617_out0) || (!v$_193_out0) && v$SUB_4617_out0);
assign v$G16_11037_out0 = ((v$_195_out0 && !v$SUB_4619_out0) || (!v$_195_out0) && v$SUB_4619_out0);
assign v$WENLS_11261_out0 = v$WENLS_601_out0;
assign v$G10_13216_out0 = ((v$_330_out0 && !v$SUB_4617_out0) || (!v$_330_out0) && v$SUB_4617_out0);
assign v$G10_13218_out0 = ((v$_332_out0 && !v$SUB_4619_out0) || (!v$_332_out0) && v$SUB_4619_out0);
assign v$G9_13286_out0 = ((v$_8749_out0 && !v$SUB_4617_out0) || (!v$_8749_out0) && v$SUB_4617_out0);
assign v$G9_13288_out0 = ((v$_8751_out0 && !v$SUB_4619_out0) || (!v$_8751_out0) && v$SUB_4619_out0);
assign v$G11_13343_out0 = ((v$_10863_out0 && !v$SUB_4617_out0) || (!v$_10863_out0) && v$SUB_4617_out0);
assign v$G11_13345_out0 = ((v$_10865_out0 && !v$SUB_4619_out0) || (!v$_10865_out0) && v$SUB_4619_out0);
assign v$G6_13638_out0 = ((v$_10378_out0 && !v$SUB_4617_out0) || (!v$_10378_out0) && v$SUB_4617_out0);
assign v$G6_13640_out0 = ((v$_10380_out0 && !v$SUB_4619_out0) || (!v$_10380_out0) && v$SUB_4619_out0);
assign v$G1_13758_out0 = ((v$_322_out0 && !v$SUB_4617_out0) || (!v$_322_out0) && v$SUB_4617_out0);
assign v$G1_13760_out0 = ((v$_324_out0 && !v$SUB_4619_out0) || (!v$_324_out0) && v$SUB_4619_out0);
assign v$WWNELS0_385_out0 = v$WENLS_11261_out0;
assign v$WEN3_1691_out0 = v$MUX6_8758_out0;
assign v$_1952_out0 = { v$G1_13758_out0,v$G2_7026_out0 };
assign v$_1954_out0 = { v$G1_13760_out0,v$G2_7028_out0 };
assign v$STALL$DUAL$CORE_1958_out0 = v$STALL$DUAL$CORE_1738_out0;
assign v$_2771_out0 = { v$SIG$RM_1767_out0,v$G2_7015_out0 };
assign v$_2772_out0 = { v$SIG$RM_1768_out0,v$G2_7016_out0 };
assign v$BYTE$READY_2853_out0 = v$BYTE$READY_10559_out0;
assign v$_4605_out0 = v$D_623_out0[0:0];
assign v$_4605_out1 = v$D_623_out0[1:1];
assign v$_4606_out0 = v$D_624_out0[0:0];
assign v$_4606_out1 = v$D_624_out0[1:1];
assign v$STALL$DUAL$CORE_4695_out0 = v$STALL$DUAL$CORE_1738_out0;
assign v$_4856_out0 = v$MUX1_31_out0[0:0];
assign v$_4856_out1 = v$MUX1_31_out0[15:15];
assign v$_4857_out0 = v$MUX1_32_out0[0:0];
assign v$_4857_out1 = v$MUX1_32_out0[15:15];
assign v$_5850_out0 = { v$_2969_out0,v$G5_230_out0 };
assign v$_7714_out0 = { v$SIG$RD_11298_out0,v$G1_646_out0 };
assign v$_7715_out0 = { v$SIG$RD_11299_out0,v$G1_647_out0 };
assign v$STALL$DUAL$CORE_12234_out0 = v$STALL$DUAL$CORE_3264_out0;
assign v$MUX13_13647_out0 = v$EQ1_2597_out0 ? v$0B00001_10554_out0 : v$RD$EXP_2601_out0;
assign v$MUX13_13648_out0 = v$EQ1_2598_out0 ? v$0B00001_10555_out0 : v$RD$EXP_2602_out0;
assign v$MUX12_13783_out0 = v$EQ2_1753_out0 ? v$0B00001_10554_out0 : v$OP2$EXP_10383_out0;
assign v$MUX12_13784_out0 = v$EQ2_1754_out0 ? v$0B00001_10555_out0 : v$OP2$EXP_10384_out0;
assign v$_97_out0 = { v$_5850_out0,v$G6_2417_out0 };
assign v$G30_183_out0 = v$G2_1887_out0 && v$STALL$DUAL$CORE_12234_out0;
assign v$G22_1899_out0 = v$G11_13439_out0 && v$STALL$DUAL$CORE_4695_out0;
assign v$NOTUSED_1968_out0 = v$_4856_out0;
assign v$NOTUSED_1969_out0 = v$_4857_out0;
assign v$SIG$RD$11bit_3301_out0 = v$_7714_out0;
assign v$SIG$RD$11bit_3302_out0 = v$_7715_out0;
assign v$SIG$RM$11bit_6892_out0 = v$_2771_out0;
assign v$SIG$RM$11bit_6893_out0 = v$_2772_out0;
assign v$STALL$dual$core_8741_out0 = v$STALL$DUAL$CORE_1958_out0;
assign v$D1_8843_out0 = (v$AD3_10483_out0 == 2'b00) ? v$WEN3_1691_out0 : 1'h0;
assign v$D1_8843_out1 = (v$AD3_10483_out0 == 2'b01) ? v$WEN3_1691_out0 : 1'h0;
assign v$D1_8843_out2 = (v$AD3_10483_out0 == 2'b10) ? v$WEN3_1691_out0 : 1'h0;
assign v$D1_8843_out3 = (v$AD3_10483_out0 == 2'b11) ? v$WEN3_1691_out0 : 1'h0;
assign v$_9805_out0 = { v$_1952_out0,v$G3_207_out0 };
assign v$_9807_out0 = { v$_1954_out0,v$G3_209_out0 };
assign v$_10262_out0 = { v$MUX13_13647_out0,v$0_10706_out0 };
assign v$_10263_out0 = { v$MUX13_13648_out0,v$0_10707_out0 };
assign v$_10370_out0 = { v$STALL$DUAL$CORE_4695_out0,v$C_1807_out0 };
assign v$_10814_out0 = { v$_4856_out1,v$C1_604_out0 };
assign v$_10815_out0 = { v$_4857_out1,v$C1_605_out0 };
assign v$_10858_out0 = { v$MUX12_13783_out0,v$0_10706_out0 };
assign v$_10859_out0 = { v$MUX12_13784_out0,v$0_10707_out0 };
assign v$OP2$SIG11_14_out0 = v$SIG$RM$11bit_6892_out0;
assign v$OP2$SIG11_15_out0 = v$SIG$RM$11bit_6893_out0;
assign v$_73_out0 = { v$_97_out0,v$G7_4822_out0 };
assign v$G4_219_out0 = v$G30_183_out0 || v$G3_2903_out0;
assign v$XOR3_2546_out0 = v$NEG1_6921_out0 ^ v$_10858_out0;
assign v$XOR3_2547_out0 = v$NEG1_6922_out0 ^ v$_10859_out0;
assign v$SUB_2909_out0 = v$G22_1899_out0;
assign v$MUX2_3255_out0 = v$LSR_6912_out0 ? v$_10814_out0 : v$MUX1_31_out0;
assign v$MUX2_3256_out0 = v$LSR_6913_out0 ? v$_10815_out0 : v$MUX1_32_out0;
assign v$EN_7093_out0 = v$STALL$dual$core_8741_out0;
assign v$_8688_out0 = { v$_9805_out0,v$G4_10998_out0 };
assign v$_8690_out0 = { v$_9807_out0,v$G4_11000_out0 };
assign v$RD$SIG11_8854_out0 = v$SIG$RD$11bit_3301_out0;
assign v$RD$SIG11_8855_out0 = v$SIG$RD$11bit_3302_out0;
assign v$A_10821_out0 = v$_10370_out0;
assign v$_60_out0 = v$A_10821_out0[10:10];
assign v$_171_out0 = v$A_10821_out0[7:7];
assign v$_179_out0 = v$A_10821_out0[3:3];
assign v$_287_out0 = v$A_10821_out0[2:2];
assign v$_1875_out0 = v$A_10821_out0[11:11];
assign v$_2022_out0 = v$A_10821_out0[5:5];
assign v$_2268_out0 = v$A_10821_out0[8:8];
assign v$_3123_out0 = v$A_10821_out0[1:1];
assign v$_3252_out0 = { v$_8688_out0,v$G5_10569_out0 };
assign v$_3254_out0 = { v$_8690_out0,v$G5_10571_out0 };
assign v$_3270_out0 = v$A_10821_out0[4:4];
assign v$MUX8_4587_out0 = v$MULTI$INSTRUCTION_13308_out0 ? v$_10858_out0 : v$XOR3_2546_out0;
assign v$MUX8_4588_out0 = v$MULTI$INSTRUCTION_13309_out0 ? v$_10859_out0 : v$XOR3_2547_out0;
assign v$OP2$SIG11_4827_out0 = v$OP2$SIG11_14_out0;
assign v$OP2$SIG11_4828_out0 = v$OP2$SIG11_15_out0;
assign v$RD$SIG11_7132_out0 = v$RD$SIG11_8854_out0;
assign v$RD$SIG11_7133_out0 = v$RD$SIG11_8855_out0;
assign v$_8682_out0 = { v$_73_out0,v$G8_2025_out0 };
assign v$Q_10339_out0 = v$OP2$SIG11_14_out0;
assign v$Q_10340_out0 = v$RD$SIG11_8854_out0;
assign v$Q_10341_out0 = v$OP2$SIG11_15_out0;
assign v$Q_10342_out0 = v$RD$SIG11_8855_out0;
assign v$_11242_out0 = v$A_10821_out0[9:9];
assign v$IN_13306_out0 = v$MUX2_3255_out0;
assign v$IN_13307_out0 = v$MUX2_3256_out0;
assign v$_13396_out0 = v$A_10821_out0[6:6];
assign v$_13562_out0 = v$A_10821_out0[0:0];
assign v$WENLDST_13755_out0 = v$G4_219_out0;
assign v$G5_229_out0 = ((v$_3270_out0 && !v$SUB_2909_out0) || (!v$_3270_out0) && v$SUB_2909_out0);
assign v$G8_2024_out0 = ((v$_171_out0 && !v$SUB_2909_out0) || (!v$_171_out0) && v$SUB_2909_out0);
assign v$G9_2332_out0 = ((v$_2268_out0 && !v$SUB_2909_out0) || (!v$_2268_out0) && v$SUB_2909_out0);
assign v$G6_2416_out0 = ((v$_2022_out0 && !v$SUB_2909_out0) || (!v$_2022_out0) && v$SUB_2909_out0);
assign v$G11_2550_out0 = ((v$_60_out0 && !v$SUB_2909_out0) || (!v$_60_out0) && v$SUB_2909_out0);
assign v$G3_2621_out0 = ((v$_287_out0 && !v$SUB_2909_out0) || (!v$_287_out0) && v$SUB_2909_out0);
assign v$G10_2632_out0 = ((v$_11242_out0 && !v$SUB_2909_out0) || (!v$_11242_out0) && v$SUB_2909_out0);
assign v$WENLDST_2682_out0 = v$WENLDST_13755_out0;
assign v$_2839_out0 = { v$_8682_out0,v$G9_2333_out0 };
assign v$_2889_out0 = v$IN_13306_out0[0:0];
assign v$_2889_out1 = v$IN_13306_out0[15:15];
assign v$_2890_out0 = v$IN_13307_out0[0:0];
assign v$_2890_out1 = v$IN_13307_out0[15:15];
assign v$G2_3239_out0 = ((v$_3123_out0 && !v$SUB_2909_out0) || (!v$_3123_out0) && v$SUB_2909_out0);
assign v$G12_4699_out0 = ((v$_1875_out0 && !v$SUB_2909_out0) || (!v$_1875_out0) && v$SUB_2909_out0);
assign v$G7_4821_out0 = ((v$_13396_out0 && !v$SUB_2909_out0) || (!v$_13396_out0) && v$SUB_2909_out0);
assign v$_7638_out0 = { v$Q_10339_out0,v$C1_10313_out0 };
assign v$_7639_out0 = { v$Q_10340_out0,v$C1_10314_out0 };
assign v$_7640_out0 = { v$Q_10341_out0,v$C1_10315_out0 };
assign v$_7641_out0 = { v$Q_10342_out0,v$C1_10316_out0 };
assign v$_10299_out0 = { v$_3252_out0,v$G6_13638_out0 };
assign v$_10301_out0 = { v$_3254_out0,v$G6_13640_out0 };
assign v$G1_10477_out0 = ((v$_13562_out0 && !v$SUB_2909_out0) || (!v$_13562_out0) && v$SUB_2909_out0);
assign v$_10808_out0 = v$IN_13306_out0[15:15];
assign v$_10809_out0 = v$IN_13307_out0[15:15];
assign v$G4_12238_out0 = ((v$_179_out0 && !v$SUB_2909_out0) || (!v$_179_out0) && v$SUB_2909_out0);
assign {v$A4_13603_out1,v$A4_13603_out0 } = v$_10262_out0 + v$MUX8_4587_out0 + v$G4_13702_out0;
assign {v$A4_13604_out1,v$A4_13604_out0 } = v$_10263_out0 + v$MUX8_4588_out0 + v$G4_13703_out0;
assign v$_120_out0 = { v$_10299_out0,v$G7_2780_out0 };
assign v$_122_out0 = { v$_10301_out0,v$G7_2782_out0 };
assign v$_333_out0 = { v$_2889_out1,v$_10808_out0 };
assign v$_334_out0 = { v$_2890_out1,v$_10809_out0 };
assign v$WENLS_600_out0 = v$WENLDST_2682_out0;
assign v$_1707_out0 = { v$G1_10477_out0,v$G2_3239_out0 };
assign v$_2650_out0 = { v$_2839_out0,v$G10_2633_out0 };
assign v$UNUSED1_3016_out0 = v$A4_13603_out1;
assign v$UNUSED1_3017_out0 = v$A4_13604_out1;
assign v$NOTUSED_4463_out0 = v$_2889_out0;
assign v$NOTUSED_4464_out0 = v$_2890_out0;
assign v$EXP$SUM_5844_out0 = v$A4_13603_out0;
assign v$EXP$SUM_5845_out0 = v$A4_13604_out0;
assign v$OUT_7708_out0 = v$_7638_out0;
assign v$OUT_7709_out0 = v$_7639_out0;
assign v$OUT_7710_out0 = v$_7640_out0;
assign v$OUT_7711_out0 = v$_7641_out0;
assign v$MUX3_8817_out0 = v$IR15_2464_out0 ? v$WENALU_8659_out0 : v$WENLDST_2682_out0;
assign v$SEL2_10323_out0 = v$A4_13603_out0[5:5];
assign v$SEL2_10324_out0 = v$A4_13604_out0[5:5];
assign v$RD$MULTI_45_out0 = v$OUT_7709_out0;
assign v$RD$MULTI_46_out0 = v$OUT_7711_out0;
assign v$RM$MULTI_210_out0 = v$OUT_7708_out0;
assign v$RM$MULTI_211_out0 = v$OUT_7710_out0;
assign v$_2386_out0 = { v$_1707_out0,v$G3_2621_out0 };
assign {v$A6_3957_out1,v$A6_3957_out0 } = v$EXP$SUM_5844_out0 + v$MUX10_10395_out0 + v$0_10706_out0;
assign {v$A6_3958_out1,v$A6_3958_out0 } = v$EXP$SUM_5845_out0 + v$MUX10_10396_out0 + v$0_10707_out0;
assign v$_4734_out0 = { v$_2650_out0,v$G11_2551_out0 };
assign v$XOR4_6960_out0 = v$EXP$SUM_5844_out0 ^ v$NEG1_6921_out0;
assign v$XOR4_6961_out0 = v$EXP$SUM_5845_out0 ^ v$NEG1_6922_out0;
assign v$MUX6_8757_out0 = v$MULTI$OPCODE_3020_out0 ? v$WEN$MULTI_2388_out0 : v$MUX3_8817_out0;
assign v$OUT_11234_out0 = v$_333_out0;
assign v$OUT_11235_out0 = v$_334_out0;
assign v$NEGATIVE_11256_out0 = v$SEL2_10323_out0;
assign v$NEGATIVE_11257_out0 = v$SEL2_10324_out0;
assign v$WENLS_11260_out0 = v$WENLS_600_out0;
assign v$_13791_out0 = { v$_120_out0,v$G8_1216_out0 };
assign v$_13793_out0 = { v$_122_out0,v$G8_1218_out0 };
assign v$WWNELS1_47_out0 = v$WENLS_11260_out0;
assign v$MUX4_275_out0 = v$NEGATIVE_11256_out0 ? v$OP2$EXP_10383_out0 : v$RD$EXP_2601_out0;
assign v$MUX4_276_out0 = v$NEGATIVE_11257_out0 ? v$OP2$EXP_10384_out0 : v$RD$EXP_2602_out0;
assign v$_465_out0 = { v$_13791_out0,v$G9_13286_out0 };
assign v$_467_out0 = { v$_13793_out0,v$G9_13288_out0 };
assign v$RM$MULTI_648_out0 = v$RM$MULTI_210_out0;
assign v$RM$MULTI_649_out0 = v$RM$MULTI_211_out0;
assign v$WEN3_1690_out0 = v$MUX6_8757_out0;
assign v$UNUSED2_2193_out0 = v$A6_3957_out1;
assign v$UNUSED2_2194_out0 = v$A6_3958_out1;
assign v$SHIFT$RD_2544_out0 = v$NEGATIVE_11256_out0;
assign v$SHIFT$RD_2545_out0 = v$NEGATIVE_11257_out0;
assign {v$A5_2638_out1,v$A5_2638_out0 } = v$XOR4_6960_out0 + v$C11_13765_out0 + v$C10_1819_out0;
assign {v$A5_2639_out1,v$A5_2639_out0 } = v$XOR4_6961_out0 + v$C11_13766_out0 + v$C10_1820_out0;
assign v$RD$FLOATING_2823_out0 = v$RD$MULTI_45_out0;
assign v$RD$FLOATING_2824_out0 = v$RD$MULTI_46_out0;
assign v$_2968_out0 = { v$_2386_out0,v$G4_12238_out0 };
assign v$SEL4_5790_out0 = v$A6_3957_out0[4:0];
assign v$SEL4_5791_out0 = v$A6_3958_out0[4:0];
assign v$MUX3_7075_out0 = v$ASR_8754_out0 ? v$OUT_11234_out0 : v$MUX2_3255_out0;
assign v$MUX3_7076_out0 = v$ASR_8755_out0 ? v$OUT_11235_out0 : v$MUX2_3256_out0;
assign v$_10784_out0 = { v$_4734_out0,v$G12_4700_out0 };
assign v$MUX11_86_out0 = v$G5_7106_out0 ? v$SEL4_5790_out0 : v$MUX4_275_out0;
assign v$MUX11_87_out0 = v$G5_7107_out0 ? v$SEL4_5791_out0 : v$MUX4_276_out0;
assign v$UNUSED_339_out0 = v$A5_2638_out1;
assign v$UNUSED_340_out0 = v$A5_2639_out1;
assign v$_423_out0 = { v$_465_out0,v$G10_13216_out0 };
assign v$_425_out0 = { v$_467_out0,v$G10_13218_out0 };
assign v$MUX7_1165_out0 = v$FLOATING$INS_13797_out0 ? v$RD$FLOATING_2823_out0 : v$RD_501_out0;
assign v$MUX7_1166_out0 = v$FLOATING$INS_13798_out0 ? v$RD$FLOATING_2824_out0 : v$RD_502_out0;
assign v$MUX8_1907_out0 = v$FLOATING$INS_13797_out0 ? v$RM$MULTI_648_out0 : v$RM_13750_out0;
assign v$MUX8_1908_out0 = v$FLOATING$INS_13798_out0 ? v$RM$MULTI_649_out0 : v$RM_13751_out0;
assign v$_2984_out0 = v$MUX3_7075_out0[0:0];
assign v$_2984_out1 = v$MUX3_7075_out0[15:15];
assign v$_2985_out0 = v$MUX3_7076_out0[0:0];
assign v$_2985_out1 = v$MUX3_7076_out0[15:15];
assign v$_5849_out0 = { v$_2968_out0,v$G5_229_out0 };
assign v$D1_8842_out0 = (v$AD3_10482_out0 == 2'b00) ? v$WEN3_1690_out0 : 1'h0;
assign v$D1_8842_out1 = (v$AD3_10482_out0 == 2'b01) ? v$WEN3_1690_out0 : 1'h0;
assign v$D1_8842_out2 = (v$AD3_10482_out0 == 2'b10) ? v$WEN3_1690_out0 : 1'h0;
assign v$D1_8842_out3 = (v$AD3_10482_out0 == 2'b11) ? v$WEN3_1690_out0 : 1'h0;
assign v$G1_10757_out0 = ! v$SHIFT$RD_2544_out0;
assign v$G1_10758_out0 = ! v$SHIFT$RD_2545_out0;
assign v$ADDER$IN_10996_out0 = v$_10784_out0;
assign v$MUX9_13486_out0 = v$NEGATIVE_11256_out0 ? v$A5_2638_out0 : v$EXP$SUM_5844_out0;
assign v$MUX9_13487_out0 = v$NEGATIVE_11257_out0 ? v$A5_2639_out0 : v$EXP$SUM_5845_out0;
assign v$_96_out0 = { v$_5849_out0,v$G6_2416_out0 };
assign v$SEL3_390_out0 = v$MUX9_13486_out0[4:0];
assign v$SEL3_391_out0 = v$MUX9_13487_out0[4:0];
assign v$RD_613_out0 = v$MUX7_1165_out0;
assign v$RD_614_out0 = v$MUX7_1166_out0;
assign v$_2835_out0 = { v$_423_out0,v$G11_13343_out0 };
assign v$_2837_out0 = { v$_425_out0,v$G11_13345_out0 };
assign v$RM_3272_out0 = v$MUX8_1907_out0;
assign v$RM_3273_out0 = v$MUX8_1908_out0;
assign v$_7120_out0 = { v$_2984_out1,v$_2984_out0 };
assign v$_7121_out0 = { v$_2985_out1,v$_2985_out0 };
assign v$SHIFT$WHICH$OP_10715_out0 = v$G1_10757_out0;
assign v$SHIFT$WHICH$OP_10716_out0 = v$G1_10758_out0;
assign v$EXP$ANS_10860_out0 = v$MUX11_86_out0;
assign v$EXP$ANS_10861_out0 = v$MUX11_87_out0;
assign v$_72_out0 = { v$_96_out0,v$G7_4821_out0 };
assign v$_437_out0 = v$RD_613_out0[2:2];
assign v$_438_out0 = v$RD_614_out0[2:2];
assign v$_2692_out0 = v$RD_613_out0[1:1];
assign v$_2693_out0 = v$RD_614_out0[1:1];
assign v$RM_2912_out0 = v$RM_3272_out0;
assign v$RM_2913_out0 = v$RM_3273_out0;
assign v$_3180_out0 = v$RD_613_out0[3:3];
assign v$_3181_out0 = v$RD_614_out0[3:3];
assign v$SHIFT$WHICH$OP_4459_out0 = v$SHIFT$WHICH$OP_10715_out0;
assign v$SHIFT$WHICH$OP_4460_out0 = v$SHIFT$WHICH$OP_10716_out0;
assign v$SHIFT$AMOUNT_4715_out0 = v$SEL3_390_out0;
assign v$SHIFT$AMOUNT_4716_out0 = v$SEL3_391_out0;
assign v$RD_4839_out0 = v$RD_613_out0;
assign v$RD_4840_out0 = v$RD_614_out0;
assign v$MUX4_7023_out0 = v$ROR_3288_out0 ? v$_7120_out0 : v$MUX3_7075_out0;
assign v$MUX4_7024_out0 = v$ROR_3289_out0 ? v$_7121_out0 : v$MUX3_7076_out0;
assign v$_7108_out0 = v$RD_613_out0[0:0];
assign v$_7109_out0 = v$RD_614_out0[0:0];
assign v$A_10274_out0 = v$RM_3272_out0;
assign v$A_10276_out0 = v$RM_3273_out0;
assign v$SHIFT$WHICH$OP_10465_out0 = v$SHIFT$WHICH$OP_10715_out0;
assign v$SHIFT$WHICH$OP_10466_out0 = v$SHIFT$WHICH$OP_10716_out0;
assign v$EXP$PRE$ANS_10765_out0 = v$EXP$ANS_10860_out0;
assign v$EXP$PRE$ANS_10766_out0 = v$EXP$ANS_10861_out0;
assign v$RM_11064_out0 = v$RM_3272_out0;
assign v$RM_11065_out0 = v$RM_3272_out0;
assign v$RM_11067_out0 = v$RM_3272_out0;
assign v$RM_11079_out0 = v$RM_3273_out0;
assign v$RM_11080_out0 = v$RM_3273_out0;
assign v$RM_11082_out0 = v$RM_3273_out0;
assign v$_11138_out0 = { v$_2835_out0,v$G12_3346_out0 };
assign v$_11140_out0 = { v$_2837_out0,v$G12_3348_out0 };
assign v$_0_out0 = v$A_10274_out0[4:4];
assign v$_2_out0 = v$A_10276_out0[4:4];
assign v$_37_out0 = v$RD_4839_out0[7:7];
assign v$_38_out0 = v$RD_4840_out0[7:7];
assign v$SHIFT$AMOUNT_226_out0 = v$SHIFT$AMOUNT_4715_out0;
assign v$SHIFT$AMOUNT_227_out0 = v$SHIFT$AMOUNT_4716_out0;
assign v$_504_out0 = v$RM_11064_out0[5:5];
assign v$_505_out0 = v$RM_11065_out0[5:5];
assign v$_507_out0 = v$RM_11067_out0[5:5];
assign v$_519_out0 = v$RM_11079_out0[5:5];
assign v$_520_out0 = v$RM_11080_out0[5:5];
assign v$_522_out0 = v$RM_11082_out0[5:5];
assign v$_569_out0 = v$RM_11064_out0[1:1];
assign v$_570_out0 = v$RM_11065_out0[1:1];
assign v$_572_out0 = v$RM_11067_out0[1:1];
assign v$_584_out0 = v$RM_11079_out0[1:1];
assign v$_585_out0 = v$RM_11080_out0[1:1];
assign v$_587_out0 = v$RM_11082_out0[1:1];
assign v$_1176_out0 = v$RD_4839_out0[13:13];
assign v$_1177_out0 = v$RD_4840_out0[13:13];
assign v$_1193_out0 = v$RD_4839_out0[4:4];
assign v$_1194_out0 = v$RD_4840_out0[4:4];
assign v$_1692_out0 = v$A_10274_out0[5:5];
assign v$_1694_out0 = v$A_10276_out0[5:5];
assign v$_1747_out0 = v$A_10274_out0[11:11];
assign v$_1749_out0 = v$A_10276_out0[11:11];
assign v$_1893_out0 = v$A_10274_out0[0:0];
assign v$_1895_out0 = v$A_10276_out0[0:0];
assign v$_1976_out0 = v$RM_11064_out0[15:15];
assign v$_1977_out0 = v$RM_11065_out0[15:15];
assign v$_1979_out0 = v$RM_11067_out0[15:15];
assign v$_1991_out0 = v$RM_11079_out0[15:15];
assign v$_1992_out0 = v$RM_11080_out0[15:15];
assign v$_1994_out0 = v$RM_11082_out0[15:15];
assign v$_2064_out0 = v$RM_11064_out0[10:10];
assign v$_2065_out0 = v$RM_11065_out0[10:10];
assign v$_2067_out0 = v$RM_11067_out0[10:10];
assign v$_2079_out0 = v$RM_11079_out0[10:10];
assign v$_2080_out0 = v$RM_11080_out0[10:10];
assign v$_2082_out0 = v$RM_11082_out0[10:10];
assign v$_2150_out0 = v$A_10274_out0[2:2];
assign v$_2152_out0 = v$A_10276_out0[2:2];
assign v$_2274_out0 = v$RM_11064_out0[12:12];
assign v$_2275_out0 = v$RM_11065_out0[12:12];
assign v$_2277_out0 = v$RM_11067_out0[12:12];
assign v$_2289_out0 = v$RM_11079_out0[12:12];
assign v$_2290_out0 = v$RM_11080_out0[12:12];
assign v$_2292_out0 = v$RM_11082_out0[12:12];
assign v$MUX1_2401_out0 = v$SHIFT$WHICH$OP_10465_out0 ? v$_2771_out0 : v$_7714_out0;
assign v$MUX1_2402_out0 = v$SHIFT$WHICH$OP_10466_out0 ? v$_2772_out0 : v$_7715_out0;
assign v$_2467_out0 = v$RD_4839_out0[8:8];
assign v$_2468_out0 = v$RD_4840_out0[8:8];
assign v$_2727_out0 = v$RM_11064_out0[2:2];
assign v$_2728_out0 = v$RM_11065_out0[2:2];
assign v$_2730_out0 = v$RM_11067_out0[2:2];
assign v$_2742_out0 = v$RM_11079_out0[2:2];
assign v$_2743_out0 = v$RM_11080_out0[2:2];
assign v$_2745_out0 = v$RM_11082_out0[2:2];
assign v$_2760_out0 = v$A_10274_out0[15:15];
assign v$_2762_out0 = v$A_10276_out0[15:15];
assign v$_2875_out0 = v$A_10274_out0[12:12];
assign v$_2877_out0 = v$A_10276_out0[12:12];
assign v$_2879_out0 = v$A_10274_out0[3:3];
assign v$_2881_out0 = v$A_10276_out0[3:3];
assign v$EXP_2907_out0 = v$EXP$PRE$ANS_10765_out0;
assign v$EXP_2908_out0 = v$EXP$PRE$ANS_10766_out0;
assign v$_2973_out0 = v$RD_4839_out0[15:15];
assign v$_2974_out0 = v$RD_4840_out0[15:15];
assign v$_2987_out0 = v$RM_11064_out0[8:8];
assign v$_2988_out0 = v$RM_11065_out0[8:8];
assign v$_2990_out0 = v$RM_11067_out0[8:8];
assign v$_3002_out0 = v$RM_11079_out0[8:8];
assign v$_3003_out0 = v$RM_11080_out0[8:8];
assign v$_3005_out0 = v$RM_11082_out0[8:8];
assign v$_3193_out0 = { v$_11138_out0,v$G13_4706_out0 };
assign v$_3195_out0 = { v$_11140_out0,v$G13_4708_out0 };
assign v$_3199_out0 = v$RD_4839_out0[10:10];
assign v$_3200_out0 = v$RD_4840_out0[10:10];
assign v$_3247_out0 = v$A_10274_out0[8:8];
assign v$_3249_out0 = v$A_10276_out0[8:8];
assign v$RDN_3349_out0 = v$_7108_out0;
assign v$RDN_3351_out0 = v$_7109_out0;
assign v$_3803_out0 = v$RD_4839_out0[12:12];
assign v$_3804_out0 = v$RD_4840_out0[12:12];
assign v$_3911_out0 = v$RM_11064_out0[11:11];
assign v$_3912_out0 = v$RM_11065_out0[11:11];
assign v$_3914_out0 = v$RM_11067_out0[11:11];
assign v$_3926_out0 = v$RM_11079_out0[11:11];
assign v$_3927_out0 = v$RM_11080_out0[11:11];
assign v$_3929_out0 = v$RM_11082_out0[11:11];
assign v$_3962_out0 = v$RM_11064_out0[9:9];
assign v$_3963_out0 = v$RM_11065_out0[9:9];
assign v$_3965_out0 = v$RM_11067_out0[9:9];
assign v$_3977_out0 = v$RM_11079_out0[9:9];
assign v$_3978_out0 = v$RM_11080_out0[9:9];
assign v$_3980_out0 = v$RM_11082_out0[9:9];
assign v$RDN_4497_out0 = v$_2692_out0;
assign v$RDN_4498_out0 = v$_437_out0;
assign v$RDN_4500_out0 = v$_3180_out0;
assign v$RDN_4512_out0 = v$_2693_out0;
assign v$RDN_4513_out0 = v$_438_out0;
assign v$RDN_4515_out0 = v$_3181_out0;
assign v$_4597_out0 = v$A_10274_out0[10:10];
assign v$_4599_out0 = v$A_10276_out0[10:10];
assign v$_4711_out0 = v$A_10274_out0[13:13];
assign v$_4713_out0 = v$A_10276_out0[13:13];
assign v$_6831_out0 = v$RM_11064_out0[14:14];
assign v$_6832_out0 = v$RM_11065_out0[14:14];
assign v$_6834_out0 = v$RM_11067_out0[14:14];
assign v$_6846_out0 = v$RM_11079_out0[14:14];
assign v$_6847_out0 = v$RM_11080_out0[14:14];
assign v$_6849_out0 = v$RM_11082_out0[14:14];
assign v$MUX5_7017_out0 = v$EN_2330_out0 ? v$MUX4_7023_out0 : v$IN_13788_out0;
assign v$MUX5_7018_out0 = v$EN_2331_out0 ? v$MUX4_7024_out0 : v$IN_13789_out0;
assign v$_8681_out0 = { v$_72_out0,v$G8_2024_out0 };
assign v$_8848_out0 = v$A_10274_out0[14:14];
assign v$_8850_out0 = v$A_10276_out0[14:14];
assign v$_10410_out0 = v$RM_11064_out0[7:7];
assign v$_10411_out0 = v$RM_11065_out0[7:7];
assign v$_10413_out0 = v$RM_11067_out0[7:7];
assign v$_10425_out0 = v$RM_11079_out0[7:7];
assign v$_10426_out0 = v$RM_11080_out0[7:7];
assign v$_10428_out0 = v$RM_11082_out0[7:7];
assign v$_10472_out0 = v$RD_4839_out0[9:9];
assign v$_10473_out0 = v$RD_4840_out0[9:9];
assign v$_10479_out0 = v$RD_4839_out0[6:6];
assign v$_10480_out0 = v$RD_4840_out0[6:6];
assign v$_10717_out0 = v$RD_4839_out0[14:14];
assign v$_10718_out0 = v$RD_4840_out0[14:14];
assign v$_10875_out0 = v$RM_11064_out0[4:4];
assign v$_10876_out0 = v$RM_11065_out0[4:4];
assign v$_10878_out0 = v$RM_11067_out0[4:4];
assign v$_10890_out0 = v$RM_11079_out0[4:4];
assign v$_10891_out0 = v$RM_11080_out0[4:4];
assign v$_10893_out0 = v$RM_11082_out0[4:4];
assign v$_11002_out0 = v$RM_11064_out0[0:0];
assign v$_11003_out0 = v$RM_11065_out0[0:0];
assign v$_11005_out0 = v$RM_11067_out0[0:0];
assign v$_11017_out0 = v$RM_11079_out0[0:0];
assign v$_11018_out0 = v$RM_11080_out0[0:0];
assign v$_11020_out0 = v$RM_11082_out0[0:0];
assign v$RM_11063_out0 = v$RM_2912_out0;
assign v$RM_11066_out0 = v$RM_2912_out0;
assign v$RM_11068_out0 = v$RM_2912_out0;
assign v$RM_11069_out0 = v$RM_2912_out0;
assign v$RM_11070_out0 = v$RM_2912_out0;
assign v$RM_11071_out0 = v$RM_2912_out0;
assign v$RM_11072_out0 = v$RM_2912_out0;
assign v$RM_11073_out0 = v$RM_2912_out0;
assign v$RM_11074_out0 = v$RM_2912_out0;
assign v$RM_11075_out0 = v$RM_2912_out0;
assign v$RM_11076_out0 = v$RM_2912_out0;
assign v$RM_11077_out0 = v$RM_2912_out0;
assign v$RM_11078_out0 = v$RM_2913_out0;
assign v$RM_11081_out0 = v$RM_2913_out0;
assign v$RM_11083_out0 = v$RM_2913_out0;
assign v$RM_11084_out0 = v$RM_2913_out0;
assign v$RM_11085_out0 = v$RM_2913_out0;
assign v$RM_11086_out0 = v$RM_2913_out0;
assign v$RM_11087_out0 = v$RM_2913_out0;
assign v$RM_11088_out0 = v$RM_2913_out0;
assign v$RM_11089_out0 = v$RM_2913_out0;
assign v$RM_11090_out0 = v$RM_2913_out0;
assign v$RM_11091_out0 = v$RM_2913_out0;
assign v$RM_11092_out0 = v$RM_2913_out0;
assign v$_11099_out0 = v$RM_11064_out0[3:3];
assign v$_11100_out0 = v$RM_11065_out0[3:3];
assign v$_11102_out0 = v$RM_11067_out0[3:3];
assign v$_11114_out0 = v$RM_11079_out0[3:3];
assign v$_11115_out0 = v$RM_11080_out0[3:3];
assign v$_11117_out0 = v$RM_11082_out0[3:3];
assign v$_11149_out0 = v$A_10274_out0[6:6];
assign v$_11151_out0 = v$A_10276_out0[6:6];
assign v$_13384_out0 = v$A_10274_out0[7:7];
assign v$_13386_out0 = v$A_10276_out0[7:7];
assign v$_13400_out0 = v$RM_11064_out0[6:6];
assign v$_13401_out0 = v$RM_11065_out0[6:6];
assign v$_13403_out0 = v$RM_11067_out0[6:6];
assign v$_13415_out0 = v$RM_11079_out0[6:6];
assign v$_13416_out0 = v$RM_11080_out0[6:6];
assign v$_13418_out0 = v$RM_11082_out0[6:6];
assign v$_13435_out0 = v$RD_4839_out0[5:5];
assign v$_13436_out0 = v$RD_4840_out0[5:5];
assign v$_13512_out0 = v$A_10274_out0[1:1];
assign v$_13514_out0 = v$A_10276_out0[1:1];
assign v$_13601_out0 = v$RD_4839_out0[11:11];
assign v$_13602_out0 = v$RD_4840_out0[11:11];
assign v$_13627_out0 = v$A_10274_out0[9:9];
assign v$_13629_out0 = v$A_10276_out0[9:9];
assign v$_13716_out0 = v$RM_11064_out0[13:13];
assign v$_13717_out0 = v$RM_11065_out0[13:13];
assign v$_13719_out0 = v$RM_11067_out0[13:13];
assign v$_13731_out0 = v$RM_11079_out0[13:13];
assign v$_13732_out0 = v$RM_11080_out0[13:13];
assign v$_13734_out0 = v$RM_11082_out0[13:13];
assign v$_174_out0 = { v$_3193_out0,v$G14_4534_out0 };
assign v$_176_out0 = { v$_3195_out0,v$G14_4536_out0 };
assign v$G3_242_out0 = v$RDN_4497_out0 && v$_2727_out0;
assign v$G3_243_out0 = v$RDN_4498_out0 && v$_2728_out0;
assign v$G3_245_out0 = v$RDN_4500_out0 && v$_2730_out0;
assign v$G3_257_out0 = v$RDN_4512_out0 && v$_2742_out0;
assign v$G3_258_out0 = v$RDN_4513_out0 && v$_2743_out0;
assign v$G3_260_out0 = v$RDN_4515_out0 && v$_2745_out0;
assign v$G4_342_out0 = v$RDN_4497_out0 && v$_11099_out0;
assign v$G4_343_out0 = v$RDN_4498_out0 && v$_11100_out0;
assign v$G4_345_out0 = v$RDN_4500_out0 && v$_11102_out0;
assign v$G4_357_out0 = v$RDN_4512_out0 && v$_11114_out0;
assign v$G4_358_out0 = v$RDN_4513_out0 && v$_11115_out0;
assign v$G4_360_out0 = v$RDN_4515_out0 && v$_11117_out0;
assign v$_503_out0 = v$RM_11063_out0[5:5];
assign v$_506_out0 = v$RM_11066_out0[5:5];
assign v$_508_out0 = v$RM_11068_out0[5:5];
assign v$_509_out0 = v$RM_11069_out0[5:5];
assign v$_510_out0 = v$RM_11070_out0[5:5];
assign v$_511_out0 = v$RM_11071_out0[5:5];
assign v$_512_out0 = v$RM_11072_out0[5:5];
assign v$_513_out0 = v$RM_11073_out0[5:5];
assign v$_514_out0 = v$RM_11074_out0[5:5];
assign v$_515_out0 = v$RM_11075_out0[5:5];
assign v$_516_out0 = v$RM_11076_out0[5:5];
assign v$_517_out0 = v$RM_11077_out0[5:5];
assign v$_518_out0 = v$RM_11078_out0[5:5];
assign v$_521_out0 = v$RM_11081_out0[5:5];
assign v$_523_out0 = v$RM_11083_out0[5:5];
assign v$_524_out0 = v$RM_11084_out0[5:5];
assign v$_525_out0 = v$RM_11085_out0[5:5];
assign v$_526_out0 = v$RM_11086_out0[5:5];
assign v$_527_out0 = v$RM_11087_out0[5:5];
assign v$_528_out0 = v$RM_11088_out0[5:5];
assign v$_529_out0 = v$RM_11089_out0[5:5];
assign v$_530_out0 = v$RM_11090_out0[5:5];
assign v$_531_out0 = v$RM_11091_out0[5:5];
assign v$_532_out0 = v$RM_11092_out0[5:5];
assign v$G8_548_out0 = v$_13384_out0 && v$RDN_3349_out0;
assign v$G8_550_out0 = v$_13386_out0 && v$RDN_3351_out0;
assign v$_568_out0 = v$RM_11063_out0[1:1];
assign v$_571_out0 = v$RM_11066_out0[1:1];
assign v$_573_out0 = v$RM_11068_out0[1:1];
assign v$_574_out0 = v$RM_11069_out0[1:1];
assign v$_575_out0 = v$RM_11070_out0[1:1];
assign v$_576_out0 = v$RM_11071_out0[1:1];
assign v$_577_out0 = v$RM_11072_out0[1:1];
assign v$_578_out0 = v$RM_11073_out0[1:1];
assign v$_579_out0 = v$RM_11074_out0[1:1];
assign v$_580_out0 = v$RM_11075_out0[1:1];
assign v$_581_out0 = v$RM_11076_out0[1:1];
assign v$_582_out0 = v$RM_11077_out0[1:1];
assign v$_583_out0 = v$RM_11078_out0[1:1];
assign v$_586_out0 = v$RM_11081_out0[1:1];
assign v$_588_out0 = v$RM_11083_out0[1:1];
assign v$_589_out0 = v$RM_11084_out0[1:1];
assign v$_590_out0 = v$RM_11085_out0[1:1];
assign v$_591_out0 = v$RM_11086_out0[1:1];
assign v$_592_out0 = v$RM_11087_out0[1:1];
assign v$_593_out0 = v$RM_11088_out0[1:1];
assign v$_594_out0 = v$RM_11089_out0[1:1];
assign v$_595_out0 = v$RM_11090_out0[1:1];
assign v$_596_out0 = v$RM_11091_out0[1:1];
assign v$_597_out0 = v$RM_11092_out0[1:1];
assign v$G14_615_out0 = v$_4711_out0 && v$RDN_3349_out0;
assign v$G14_617_out0 = v$_4713_out0 && v$RDN_3351_out0;
assign v$G13_642_out0 = v$_2875_out0 && v$RDN_3349_out0;
assign v$G13_644_out0 = v$_2877_out0 && v$RDN_3351_out0;
assign v$OUT_1136_out0 = v$MUX5_7017_out0;
assign v$OUT_1137_out0 = v$MUX5_7018_out0;
assign v$G2_1809_out0 = v$_13512_out0 && v$RDN_3349_out0;
assign v$G2_1811_out0 = v$_13514_out0 && v$RDN_3351_out0;
assign v$G1_1879_out0 = v$_1893_out0 && v$RDN_3349_out0;
assign v$G1_1881_out0 = v$_1895_out0 && v$RDN_3351_out0;
assign v$G1_1910_out0 = v$RDN_4497_out0 && v$_569_out0;
assign v$G1_1911_out0 = v$RDN_4498_out0 && v$_570_out0;
assign v$G1_1913_out0 = v$RDN_4500_out0 && v$_572_out0;
assign v$G1_1925_out0 = v$RDN_4512_out0 && v$_584_out0;
assign v$G1_1926_out0 = v$RDN_4513_out0 && v$_585_out0;
assign v$G1_1928_out0 = v$RDN_4515_out0 && v$_587_out0;
assign v$_1975_out0 = v$RM_11063_out0[15:15];
assign v$_1978_out0 = v$RM_11066_out0[15:15];
assign v$_1980_out0 = v$RM_11068_out0[15:15];
assign v$_1981_out0 = v$RM_11069_out0[15:15];
assign v$_1982_out0 = v$RM_11070_out0[15:15];
assign v$_1983_out0 = v$RM_11071_out0[15:15];
assign v$_1984_out0 = v$RM_11072_out0[15:15];
assign v$_1985_out0 = v$RM_11073_out0[15:15];
assign v$_1986_out0 = v$RM_11074_out0[15:15];
assign v$_1987_out0 = v$RM_11075_out0[15:15];
assign v$_1988_out0 = v$RM_11076_out0[15:15];
assign v$_1989_out0 = v$RM_11077_out0[15:15];
assign v$_1990_out0 = v$RM_11078_out0[15:15];
assign v$_1993_out0 = v$RM_11081_out0[15:15];
assign v$_1995_out0 = v$RM_11083_out0[15:15];
assign v$_1996_out0 = v$RM_11084_out0[15:15];
assign v$_1997_out0 = v$RM_11085_out0[15:15];
assign v$_1998_out0 = v$RM_11086_out0[15:15];
assign v$_1999_out0 = v$RM_11087_out0[15:15];
assign v$_2000_out0 = v$RM_11088_out0[15:15];
assign v$_2001_out0 = v$RM_11089_out0[15:15];
assign v$_2002_out0 = v$RM_11090_out0[15:15];
assign v$_2003_out0 = v$RM_11091_out0[15:15];
assign v$_2004_out0 = v$RM_11092_out0[15:15];
assign v$_2063_out0 = v$RM_11063_out0[10:10];
assign v$_2066_out0 = v$RM_11066_out0[10:10];
assign v$_2068_out0 = v$RM_11068_out0[10:10];
assign v$_2069_out0 = v$RM_11069_out0[10:10];
assign v$_2070_out0 = v$RM_11070_out0[10:10];
assign v$_2071_out0 = v$RM_11071_out0[10:10];
assign v$_2072_out0 = v$RM_11072_out0[10:10];
assign v$_2073_out0 = v$RM_11073_out0[10:10];
assign v$_2074_out0 = v$RM_11074_out0[10:10];
assign v$_2075_out0 = v$RM_11075_out0[10:10];
assign v$_2076_out0 = v$RM_11076_out0[10:10];
assign v$_2077_out0 = v$RM_11077_out0[10:10];
assign v$_2078_out0 = v$RM_11078_out0[10:10];
assign v$_2081_out0 = v$RM_11081_out0[10:10];
assign v$_2083_out0 = v$RM_11083_out0[10:10];
assign v$_2084_out0 = v$RM_11084_out0[10:10];
assign v$_2085_out0 = v$RM_11085_out0[10:10];
assign v$_2086_out0 = v$RM_11086_out0[10:10];
assign v$_2087_out0 = v$RM_11087_out0[10:10];
assign v$_2088_out0 = v$RM_11088_out0[10:10];
assign v$_2089_out0 = v$RM_11089_out0[10:10];
assign v$_2090_out0 = v$RM_11090_out0[10:10];
assign v$_2091_out0 = v$RM_11091_out0[10:10];
assign v$_2092_out0 = v$RM_11092_out0[10:10];
assign v$G6_2117_out0 = v$RDN_4497_out0 && v$_13400_out0;
assign v$G6_2118_out0 = v$RDN_4498_out0 && v$_13401_out0;
assign v$G6_2120_out0 = v$RDN_4500_out0 && v$_13403_out0;
assign v$G6_2132_out0 = v$RDN_4512_out0 && v$_13415_out0;
assign v$G6_2133_out0 = v$RDN_4513_out0 && v$_13416_out0;
assign v$G6_2135_out0 = v$RDN_4515_out0 && v$_13418_out0;
assign v$_2273_out0 = v$RM_11063_out0[12:12];
assign v$_2276_out0 = v$RM_11066_out0[12:12];
assign v$_2278_out0 = v$RM_11068_out0[12:12];
assign v$_2279_out0 = v$RM_11069_out0[12:12];
assign v$_2280_out0 = v$RM_11070_out0[12:12];
assign v$_2281_out0 = v$RM_11071_out0[12:12];
assign v$_2282_out0 = v$RM_11072_out0[12:12];
assign v$_2283_out0 = v$RM_11073_out0[12:12];
assign v$_2284_out0 = v$RM_11074_out0[12:12];
assign v$_2285_out0 = v$RM_11075_out0[12:12];
assign v$_2286_out0 = v$RM_11076_out0[12:12];
assign v$_2287_out0 = v$RM_11077_out0[12:12];
assign v$_2288_out0 = v$RM_11078_out0[12:12];
assign v$_2291_out0 = v$RM_11081_out0[12:12];
assign v$_2293_out0 = v$RM_11083_out0[12:12];
assign v$_2294_out0 = v$RM_11084_out0[12:12];
assign v$_2295_out0 = v$RM_11085_out0[12:12];
assign v$_2296_out0 = v$RM_11086_out0[12:12];
assign v$_2297_out0 = v$RM_11087_out0[12:12];
assign v$_2298_out0 = v$RM_11088_out0[12:12];
assign v$_2299_out0 = v$RM_11089_out0[12:12];
assign v$_2300_out0 = v$RM_11090_out0[12:12];
assign v$_2301_out0 = v$RM_11091_out0[12:12];
assign v$_2302_out0 = v$RM_11092_out0[12:12];
assign v$EXP_2441_out0 = v$EXP_2907_out0;
assign v$EXP_2442_out0 = v$EXP_2908_out0;
assign v$G8_2473_out0 = v$RDN_4497_out0 && v$_2987_out0;
assign v$G8_2474_out0 = v$RDN_4498_out0 && v$_2988_out0;
assign v$G8_2476_out0 = v$RDN_4500_out0 && v$_2990_out0;
assign v$G8_2488_out0 = v$RDN_4512_out0 && v$_3002_out0;
assign v$G8_2489_out0 = v$RDN_4513_out0 && v$_3003_out0;
assign v$G8_2491_out0 = v$RDN_4515_out0 && v$_3005_out0;
assign v$G10_2640_out0 = v$_13627_out0 && v$RDN_3349_out0;
assign v$G10_2642_out0 = v$_13629_out0 && v$RDN_3351_out0;
assign v$_2726_out0 = v$RM_11063_out0[2:2];
assign v$_2729_out0 = v$RM_11066_out0[2:2];
assign v$_2731_out0 = v$RM_11068_out0[2:2];
assign v$_2732_out0 = v$RM_11069_out0[2:2];
assign v$_2733_out0 = v$RM_11070_out0[2:2];
assign v$_2734_out0 = v$RM_11071_out0[2:2];
assign v$_2735_out0 = v$RM_11072_out0[2:2];
assign v$_2736_out0 = v$RM_11073_out0[2:2];
assign v$_2737_out0 = v$RM_11074_out0[2:2];
assign v$_2738_out0 = v$RM_11075_out0[2:2];
assign v$_2739_out0 = v$RM_11076_out0[2:2];
assign v$_2740_out0 = v$RM_11077_out0[2:2];
assign v$_2741_out0 = v$RM_11078_out0[2:2];
assign v$_2744_out0 = v$RM_11081_out0[2:2];
assign v$_2746_out0 = v$RM_11083_out0[2:2];
assign v$_2747_out0 = v$RM_11084_out0[2:2];
assign v$_2748_out0 = v$RM_11085_out0[2:2];
assign v$_2749_out0 = v$RM_11086_out0[2:2];
assign v$_2750_out0 = v$RM_11087_out0[2:2];
assign v$_2751_out0 = v$RM_11088_out0[2:2];
assign v$_2752_out0 = v$RM_11089_out0[2:2];
assign v$_2753_out0 = v$RM_11090_out0[2:2];
assign v$_2754_out0 = v$RM_11091_out0[2:2];
assign v$_2755_out0 = v$RM_11092_out0[2:2];
assign v$G4_2767_out0 = v$_2879_out0 && v$RDN_3349_out0;
assign v$G4_2769_out0 = v$_2881_out0 && v$RDN_3351_out0;
assign v$G5_2783_out0 = v$_0_out0 && v$RDN_3349_out0;
assign v$G5_2785_out0 = v$_2_out0 && v$RDN_3351_out0;
assign v$_2838_out0 = { v$_8681_out0,v$G9_2332_out0 };
assign v$G9_2895_out0 = v$_3247_out0 && v$RDN_3349_out0;
assign v$G9_2897_out0 = v$_3249_out0 && v$RDN_3351_out0;
assign v$G11_2937_out0 = v$_4597_out0 && v$RDN_3349_out0;
assign v$G11_2939_out0 = v$_4599_out0 && v$RDN_3351_out0;
assign v$_2986_out0 = v$RM_11063_out0[8:8];
assign v$_2989_out0 = v$RM_11066_out0[8:8];
assign v$_2991_out0 = v$RM_11068_out0[8:8];
assign v$_2992_out0 = v$RM_11069_out0[8:8];
assign v$_2993_out0 = v$RM_11070_out0[8:8];
assign v$_2994_out0 = v$RM_11071_out0[8:8];
assign v$_2995_out0 = v$RM_11072_out0[8:8];
assign v$_2996_out0 = v$RM_11073_out0[8:8];
assign v$_2997_out0 = v$RM_11074_out0[8:8];
assign v$_2998_out0 = v$RM_11075_out0[8:8];
assign v$_2999_out0 = v$RM_11076_out0[8:8];
assign v$_3000_out0 = v$RM_11077_out0[8:8];
assign v$_3001_out0 = v$RM_11078_out0[8:8];
assign v$_3004_out0 = v$RM_11081_out0[8:8];
assign v$_3006_out0 = v$RM_11083_out0[8:8];
assign v$_3007_out0 = v$RM_11084_out0[8:8];
assign v$_3008_out0 = v$RM_11085_out0[8:8];
assign v$_3009_out0 = v$RM_11086_out0[8:8];
assign v$_3010_out0 = v$RM_11087_out0[8:8];
assign v$_3011_out0 = v$RM_11088_out0[8:8];
assign v$_3012_out0 = v$RM_11089_out0[8:8];
assign v$_3013_out0 = v$RM_11090_out0[8:8];
assign v$_3014_out0 = v$RM_11091_out0[8:8];
assign v$_3015_out0 = v$RM_11092_out0[8:8];
assign v$_3910_out0 = v$RM_11063_out0[11:11];
assign v$_3913_out0 = v$RM_11066_out0[11:11];
assign v$_3915_out0 = v$RM_11068_out0[11:11];
assign v$_3916_out0 = v$RM_11069_out0[11:11];
assign v$_3917_out0 = v$RM_11070_out0[11:11];
assign v$_3918_out0 = v$RM_11071_out0[11:11];
assign v$_3919_out0 = v$RM_11072_out0[11:11];
assign v$_3920_out0 = v$RM_11073_out0[11:11];
assign v$_3921_out0 = v$RM_11074_out0[11:11];
assign v$_3922_out0 = v$RM_11075_out0[11:11];
assign v$_3923_out0 = v$RM_11076_out0[11:11];
assign v$_3924_out0 = v$RM_11077_out0[11:11];
assign v$_3925_out0 = v$RM_11078_out0[11:11];
assign v$_3928_out0 = v$RM_11081_out0[11:11];
assign v$_3930_out0 = v$RM_11083_out0[11:11];
assign v$_3931_out0 = v$RM_11084_out0[11:11];
assign v$_3932_out0 = v$RM_11085_out0[11:11];
assign v$_3933_out0 = v$RM_11086_out0[11:11];
assign v$_3934_out0 = v$RM_11087_out0[11:11];
assign v$_3935_out0 = v$RM_11088_out0[11:11];
assign v$_3936_out0 = v$RM_11089_out0[11:11];
assign v$_3937_out0 = v$RM_11090_out0[11:11];
assign v$_3938_out0 = v$RM_11091_out0[11:11];
assign v$_3939_out0 = v$RM_11092_out0[11:11];
assign v$B_3946_out0 = v$SHIFT$AMOUNT_226_out0;
assign v$B_3947_out0 = v$SHIFT$AMOUNT_227_out0;
assign v$_3961_out0 = v$RM_11063_out0[9:9];
assign v$_3964_out0 = v$RM_11066_out0[9:9];
assign v$_3966_out0 = v$RM_11068_out0[9:9];
assign v$_3967_out0 = v$RM_11069_out0[9:9];
assign v$_3968_out0 = v$RM_11070_out0[9:9];
assign v$_3969_out0 = v$RM_11071_out0[9:9];
assign v$_3970_out0 = v$RM_11072_out0[9:9];
assign v$_3971_out0 = v$RM_11073_out0[9:9];
assign v$_3972_out0 = v$RM_11074_out0[9:9];
assign v$_3973_out0 = v$RM_11075_out0[9:9];
assign v$_3974_out0 = v$RM_11076_out0[9:9];
assign v$_3975_out0 = v$RM_11077_out0[9:9];
assign v$_3976_out0 = v$RM_11078_out0[9:9];
assign v$_3979_out0 = v$RM_11081_out0[9:9];
assign v$_3981_out0 = v$RM_11083_out0[9:9];
assign v$_3982_out0 = v$RM_11084_out0[9:9];
assign v$_3983_out0 = v$RM_11085_out0[9:9];
assign v$_3984_out0 = v$RM_11086_out0[9:9];
assign v$_3985_out0 = v$RM_11087_out0[9:9];
assign v$_3986_out0 = v$RM_11088_out0[9:9];
assign v$_3987_out0 = v$RM_11089_out0[9:9];
assign v$_3988_out0 = v$RM_11090_out0[9:9];
assign v$_3989_out0 = v$RM_11091_out0[9:9];
assign v$_3990_out0 = v$RM_11092_out0[9:9];
assign v$RDN_4496_out0 = v$_1193_out0;
assign v$RDN_4499_out0 = v$_13601_out0;
assign v$RDN_4501_out0 = v$_3199_out0;
assign v$RDN_4502_out0 = v$_2973_out0;
assign v$RDN_4503_out0 = v$_10717_out0;
assign v$RDN_4504_out0 = v$_3803_out0;
assign v$RDN_4505_out0 = v$_2467_out0;
assign v$RDN_4506_out0 = v$_13435_out0;
assign v$RDN_4507_out0 = v$_37_out0;
assign v$RDN_4508_out0 = v$_1176_out0;
assign v$RDN_4509_out0 = v$_10479_out0;
assign v$RDN_4510_out0 = v$_10472_out0;
assign v$RDN_4511_out0 = v$_1194_out0;
assign v$RDN_4514_out0 = v$_13602_out0;
assign v$RDN_4516_out0 = v$_3200_out0;
assign v$RDN_4517_out0 = v$_2974_out0;
assign v$RDN_4518_out0 = v$_10718_out0;
assign v$RDN_4519_out0 = v$_3804_out0;
assign v$RDN_4520_out0 = v$_2468_out0;
assign v$RDN_4521_out0 = v$_13436_out0;
assign v$RDN_4522_out0 = v$_38_out0;
assign v$RDN_4523_out0 = v$_1177_out0;
assign v$RDN_4524_out0 = v$_10480_out0;
assign v$RDN_4525_out0 = v$_10473_out0;
assign v$G2_4621_out0 = v$RDN_4497_out0 && v$_10875_out0;
assign v$G2_4622_out0 = v$RDN_4498_out0 && v$_10876_out0;
assign v$G2_4624_out0 = v$RDN_4500_out0 && v$_10878_out0;
assign v$G2_4636_out0 = v$RDN_4512_out0 && v$_10890_out0;
assign v$G2_4637_out0 = v$RDN_4513_out0 && v$_10891_out0;
assign v$G2_4639_out0 = v$RDN_4515_out0 && v$_10893_out0;
assign v$G15_4654_out0 = v$_8848_out0 && v$RDN_3349_out0;
assign v$G15_4656_out0 = v$_8850_out0 && v$RDN_3351_out0;
assign v$_6830_out0 = v$RM_11063_out0[14:14];
assign v$_6833_out0 = v$RM_11066_out0[14:14];
assign v$_6835_out0 = v$RM_11068_out0[14:14];
assign v$_6836_out0 = v$RM_11069_out0[14:14];
assign v$_6837_out0 = v$RM_11070_out0[14:14];
assign v$_6838_out0 = v$RM_11071_out0[14:14];
assign v$_6839_out0 = v$RM_11072_out0[14:14];
assign v$_6840_out0 = v$RM_11073_out0[14:14];
assign v$_6841_out0 = v$RM_11074_out0[14:14];
assign v$_6842_out0 = v$RM_11075_out0[14:14];
assign v$_6843_out0 = v$RM_11076_out0[14:14];
assign v$_6844_out0 = v$RM_11077_out0[14:14];
assign v$_6845_out0 = v$RM_11078_out0[14:14];
assign v$_6848_out0 = v$RM_11081_out0[14:14];
assign v$_6850_out0 = v$RM_11083_out0[14:14];
assign v$_6851_out0 = v$RM_11084_out0[14:14];
assign v$_6852_out0 = v$RM_11085_out0[14:14];
assign v$_6853_out0 = v$RM_11086_out0[14:14];
assign v$_6854_out0 = v$RM_11087_out0[14:14];
assign v$_6855_out0 = v$RM_11088_out0[14:14];
assign v$_6856_out0 = v$RM_11089_out0[14:14];
assign v$_6857_out0 = v$RM_11090_out0[14:14];
assign v$_6858_out0 = v$RM_11091_out0[14:14];
assign v$_6859_out0 = v$RM_11092_out0[14:14];
assign v$EQ1_6956_out0 = v$EXP_2907_out0 == 5'h0;
assign v$EQ1_6957_out0 = v$EXP_2908_out0 == 5'h0;
assign v$G3_7087_out0 = v$_2150_out0 && v$RDN_3349_out0;
assign v$G3_7089_out0 = v$_2152_out0 && v$RDN_3351_out0;
assign v$G7_8655_out0 = v$_11149_out0 && v$RDN_3349_out0;
assign v$G7_8657_out0 = v$_11151_out0 && v$RDN_3351_out0;
assign v$G6_8834_out0 = v$_1692_out0 && v$RDN_3349_out0;
assign v$G6_8836_out0 = v$_1694_out0 && v$RDN_3351_out0;
assign v$_10409_out0 = v$RM_11063_out0[7:7];
assign v$_10412_out0 = v$RM_11066_out0[7:7];
assign v$_10414_out0 = v$RM_11068_out0[7:7];
assign v$_10415_out0 = v$RM_11069_out0[7:7];
assign v$_10416_out0 = v$RM_11070_out0[7:7];
assign v$_10417_out0 = v$RM_11071_out0[7:7];
assign v$_10418_out0 = v$RM_11072_out0[7:7];
assign v$_10419_out0 = v$RM_11073_out0[7:7];
assign v$_10420_out0 = v$RM_11074_out0[7:7];
assign v$_10421_out0 = v$RM_11075_out0[7:7];
assign v$_10422_out0 = v$RM_11076_out0[7:7];
assign v$_10423_out0 = v$RM_11077_out0[7:7];
assign v$_10424_out0 = v$RM_11078_out0[7:7];
assign v$_10427_out0 = v$RM_11081_out0[7:7];
assign v$_10429_out0 = v$RM_11083_out0[7:7];
assign v$_10430_out0 = v$RM_11084_out0[7:7];
assign v$_10431_out0 = v$RM_11085_out0[7:7];
assign v$_10432_out0 = v$RM_11086_out0[7:7];
assign v$_10433_out0 = v$RM_11087_out0[7:7];
assign v$_10434_out0 = v$RM_11088_out0[7:7];
assign v$_10435_out0 = v$RM_11089_out0[7:7];
assign v$_10436_out0 = v$RM_11090_out0[7:7];
assign v$_10437_out0 = v$RM_11091_out0[7:7];
assign v$_10438_out0 = v$RM_11092_out0[7:7];
assign v$G9_10573_out0 = v$RDN_4497_out0 && v$_3962_out0;
assign v$G9_10574_out0 = v$RDN_4498_out0 && v$_3963_out0;
assign v$G9_10576_out0 = v$RDN_4500_out0 && v$_3965_out0;
assign v$G9_10588_out0 = v$RDN_4512_out0 && v$_3977_out0;
assign v$G9_10589_out0 = v$RDN_4513_out0 && v$_3978_out0;
assign v$G9_10591_out0 = v$RDN_4515_out0 && v$_3980_out0;
assign v$G5_10622_out0 = v$RDN_4497_out0 && v$_504_out0;
assign v$G5_10623_out0 = v$RDN_4498_out0 && v$_505_out0;
assign v$G5_10625_out0 = v$RDN_4500_out0 && v$_507_out0;
assign v$G5_10637_out0 = v$RDN_4512_out0 && v$_519_out0;
assign v$G5_10638_out0 = v$RDN_4513_out0 && v$_520_out0;
assign v$G5_10640_out0 = v$RDN_4515_out0 && v$_522_out0;
assign v$G12_10688_out0 = v$_1747_out0 && v$RDN_3349_out0;
assign v$G12_10690_out0 = v$_1749_out0 && v$RDN_3351_out0;
assign v$SIG$TO$SHIFT_10712_out0 = v$MUX1_2401_out0;
assign v$SIG$TO$SHIFT_10713_out0 = v$MUX1_2402_out0;
assign v$_10874_out0 = v$RM_11063_out0[4:4];
assign v$_10877_out0 = v$RM_11066_out0[4:4];
assign v$_10879_out0 = v$RM_11068_out0[4:4];
assign v$_10880_out0 = v$RM_11069_out0[4:4];
assign v$_10881_out0 = v$RM_11070_out0[4:4];
assign v$_10882_out0 = v$RM_11071_out0[4:4];
assign v$_10883_out0 = v$RM_11072_out0[4:4];
assign v$_10884_out0 = v$RM_11073_out0[4:4];
assign v$_10885_out0 = v$RM_11074_out0[4:4];
assign v$_10886_out0 = v$RM_11075_out0[4:4];
assign v$_10887_out0 = v$RM_11076_out0[4:4];
assign v$_10888_out0 = v$RM_11077_out0[4:4];
assign v$_10889_out0 = v$RM_11078_out0[4:4];
assign v$_10892_out0 = v$RM_11081_out0[4:4];
assign v$_10894_out0 = v$RM_11083_out0[4:4];
assign v$_10895_out0 = v$RM_11084_out0[4:4];
assign v$_10896_out0 = v$RM_11085_out0[4:4];
assign v$_10897_out0 = v$RM_11086_out0[4:4];
assign v$_10898_out0 = v$RM_11087_out0[4:4];
assign v$_10899_out0 = v$RM_11088_out0[4:4];
assign v$_10900_out0 = v$RM_11089_out0[4:4];
assign v$_10901_out0 = v$RM_11090_out0[4:4];
assign v$_10902_out0 = v$RM_11091_out0[4:4];
assign v$_10903_out0 = v$RM_11092_out0[4:4];
assign v$G16_10906_out0 = v$_2760_out0 && v$RDN_3349_out0;
assign v$G16_10908_out0 = v$_2762_out0 && v$RDN_3351_out0;
assign v$_11001_out0 = v$RM_11063_out0[0:0];
assign v$_11004_out0 = v$RM_11066_out0[0:0];
assign v$_11006_out0 = v$RM_11068_out0[0:0];
assign v$_11007_out0 = v$RM_11069_out0[0:0];
assign v$_11008_out0 = v$RM_11070_out0[0:0];
assign v$_11009_out0 = v$RM_11071_out0[0:0];
assign v$_11010_out0 = v$RM_11072_out0[0:0];
assign v$_11011_out0 = v$RM_11073_out0[0:0];
assign v$_11012_out0 = v$RM_11074_out0[0:0];
assign v$_11013_out0 = v$RM_11075_out0[0:0];
assign v$_11014_out0 = v$RM_11076_out0[0:0];
assign v$_11015_out0 = v$RM_11077_out0[0:0];
assign v$_11016_out0 = v$RM_11078_out0[0:0];
assign v$_11019_out0 = v$RM_11081_out0[0:0];
assign v$_11021_out0 = v$RM_11083_out0[0:0];
assign v$_11022_out0 = v$RM_11084_out0[0:0];
assign v$_11023_out0 = v$RM_11085_out0[0:0];
assign v$_11024_out0 = v$RM_11086_out0[0:0];
assign v$_11025_out0 = v$RM_11087_out0[0:0];
assign v$_11026_out0 = v$RM_11088_out0[0:0];
assign v$_11027_out0 = v$RM_11089_out0[0:0];
assign v$_11028_out0 = v$RM_11090_out0[0:0];
assign v$_11029_out0 = v$RM_11091_out0[0:0];
assign v$_11030_out0 = v$RM_11092_out0[0:0];
assign v$_11098_out0 = v$RM_11063_out0[3:3];
assign v$_11101_out0 = v$RM_11066_out0[3:3];
assign v$_11103_out0 = v$RM_11068_out0[3:3];
assign v$_11104_out0 = v$RM_11069_out0[3:3];
assign v$_11105_out0 = v$RM_11070_out0[3:3];
assign v$_11106_out0 = v$RM_11071_out0[3:3];
assign v$_11107_out0 = v$RM_11072_out0[3:3];
assign v$_11108_out0 = v$RM_11073_out0[3:3];
assign v$_11109_out0 = v$RM_11074_out0[3:3];
assign v$_11110_out0 = v$RM_11075_out0[3:3];
assign v$_11111_out0 = v$RM_11076_out0[3:3];
assign v$_11112_out0 = v$RM_11077_out0[3:3];
assign v$_11113_out0 = v$RM_11078_out0[3:3];
assign v$_11116_out0 = v$RM_11081_out0[3:3];
assign v$_11118_out0 = v$RM_11083_out0[3:3];
assign v$_11119_out0 = v$RM_11084_out0[3:3];
assign v$_11120_out0 = v$RM_11085_out0[3:3];
assign v$_11121_out0 = v$RM_11086_out0[3:3];
assign v$_11122_out0 = v$RM_11087_out0[3:3];
assign v$_11123_out0 = v$RM_11088_out0[3:3];
assign v$_11124_out0 = v$RM_11089_out0[3:3];
assign v$_11125_out0 = v$RM_11090_out0[3:3];
assign v$_11126_out0 = v$RM_11091_out0[3:3];
assign v$_11127_out0 = v$RM_11092_out0[3:3];
assign v$EQ2_11254_out0 = v$EXP_2907_out0 == 5'h1;
assign v$EQ2_11255_out0 = v$EXP_2908_out0 == 5'h1;
assign v$G7_11263_out0 = v$RDN_4497_out0 && v$_10410_out0;
assign v$G7_11264_out0 = v$RDN_4498_out0 && v$_10411_out0;
assign v$G7_11266_out0 = v$RDN_4500_out0 && v$_10413_out0;
assign v$G7_11278_out0 = v$RDN_4512_out0 && v$_10425_out0;
assign v$G7_11279_out0 = v$RDN_4513_out0 && v$_10426_out0;
assign v$G7_11281_out0 = v$RDN_4515_out0 && v$_10428_out0;
assign v$G16_13184_out0 = v$RDN_4497_out0 && v$_11002_out0;
assign v$G16_13185_out0 = v$RDN_4498_out0 && v$_11003_out0;
assign v$G16_13187_out0 = v$RDN_4500_out0 && v$_11005_out0;
assign v$G16_13199_out0 = v$RDN_4512_out0 && v$_11017_out0;
assign v$G16_13200_out0 = v$RDN_4513_out0 && v$_11018_out0;
assign v$G16_13202_out0 = v$RDN_4515_out0 && v$_11020_out0;
assign v$_13399_out0 = v$RM_11063_out0[6:6];
assign v$_13402_out0 = v$RM_11066_out0[6:6];
assign v$_13404_out0 = v$RM_11068_out0[6:6];
assign v$_13405_out0 = v$RM_11069_out0[6:6];
assign v$_13406_out0 = v$RM_11070_out0[6:6];
assign v$_13407_out0 = v$RM_11071_out0[6:6];
assign v$_13408_out0 = v$RM_11072_out0[6:6];
assign v$_13409_out0 = v$RM_11073_out0[6:6];
assign v$_13410_out0 = v$RM_11074_out0[6:6];
assign v$_13411_out0 = v$RM_11075_out0[6:6];
assign v$_13412_out0 = v$RM_11076_out0[6:6];
assign v$_13413_out0 = v$RM_11077_out0[6:6];
assign v$_13414_out0 = v$RM_11078_out0[6:6];
assign v$_13417_out0 = v$RM_11081_out0[6:6];
assign v$_13419_out0 = v$RM_11083_out0[6:6];
assign v$_13420_out0 = v$RM_11084_out0[6:6];
assign v$_13421_out0 = v$RM_11085_out0[6:6];
assign v$_13422_out0 = v$RM_11086_out0[6:6];
assign v$_13423_out0 = v$RM_11087_out0[6:6];
assign v$_13424_out0 = v$RM_11088_out0[6:6];
assign v$_13425_out0 = v$RM_11089_out0[6:6];
assign v$_13426_out0 = v$RM_11090_out0[6:6];
assign v$_13427_out0 = v$RM_11091_out0[6:6];
assign v$_13428_out0 = v$RM_11092_out0[6:6];
assign v$RD_13568_out0 = v$RDN_4497_out0;
assign v$RD_13569_out0 = v$RDN_4498_out0;
assign v$RD_13571_out0 = v$RDN_4500_out0;
assign v$RD_13583_out0 = v$RDN_4512_out0;
assign v$RD_13584_out0 = v$RDN_4513_out0;
assign v$RD_13586_out0 = v$RDN_4515_out0;
assign v$_13715_out0 = v$RM_11063_out0[13:13];
assign v$_13718_out0 = v$RM_11066_out0[13:13];
assign v$_13720_out0 = v$RM_11068_out0[13:13];
assign v$_13721_out0 = v$RM_11069_out0[13:13];
assign v$_13722_out0 = v$RM_11070_out0[13:13];
assign v$_13723_out0 = v$RM_11071_out0[13:13];
assign v$_13724_out0 = v$RM_11072_out0[13:13];
assign v$_13725_out0 = v$RM_11073_out0[13:13];
assign v$_13726_out0 = v$RM_11074_out0[13:13];
assign v$_13727_out0 = v$RM_11075_out0[13:13];
assign v$_13728_out0 = v$RM_11076_out0[13:13];
assign v$_13729_out0 = v$RM_11077_out0[13:13];
assign v$_13730_out0 = v$RM_11078_out0[13:13];
assign v$_13733_out0 = v$RM_11081_out0[13:13];
assign v$_13735_out0 = v$RM_11083_out0[13:13];
assign v$_13736_out0 = v$RM_11084_out0[13:13];
assign v$_13737_out0 = v$RM_11085_out0[13:13];
assign v$_13738_out0 = v$RM_11086_out0[13:13];
assign v$_13739_out0 = v$RM_11087_out0[13:13];
assign v$_13740_out0 = v$RM_11088_out0[13:13];
assign v$_13741_out0 = v$RM_11089_out0[13:13];
assign v$_13742_out0 = v$RM_11090_out0[13:13];
assign v$_13743_out0 = v$RM_11091_out0[13:13];
assign v$_13744_out0 = v$RM_11092_out0[13:13];
assign v$G15_133_out0 = v$RD_13568_out0 && v$_1976_out0;
assign v$G15_134_out0 = v$RD_13569_out0 && v$_1977_out0;
assign v$G15_136_out0 = v$RD_13571_out0 && v$_1979_out0;
assign v$G15_148_out0 = v$RD_13583_out0 && v$_1991_out0;
assign v$G15_149_out0 = v$RD_13584_out0 && v$_1992_out0;
assign v$G15_151_out0 = v$RD_13586_out0 && v$_1994_out0;
assign v$G3_241_out0 = v$RDN_4496_out0 && v$_2726_out0;
assign v$G3_244_out0 = v$RDN_4499_out0 && v$_2729_out0;
assign v$G3_246_out0 = v$RDN_4501_out0 && v$_2731_out0;
assign v$G3_247_out0 = v$RDN_4502_out0 && v$_2732_out0;
assign v$G3_248_out0 = v$RDN_4503_out0 && v$_2733_out0;
assign v$G3_249_out0 = v$RDN_4504_out0 && v$_2734_out0;
assign v$G3_250_out0 = v$RDN_4505_out0 && v$_2735_out0;
assign v$G3_251_out0 = v$RDN_4506_out0 && v$_2736_out0;
assign v$G3_252_out0 = v$RDN_4507_out0 && v$_2737_out0;
assign v$G3_253_out0 = v$RDN_4508_out0 && v$_2738_out0;
assign v$G3_254_out0 = v$RDN_4509_out0 && v$_2739_out0;
assign v$G3_255_out0 = v$RDN_4510_out0 && v$_2740_out0;
assign v$G3_256_out0 = v$RDN_4511_out0 && v$_2741_out0;
assign v$G3_259_out0 = v$RDN_4514_out0 && v$_2744_out0;
assign v$G3_261_out0 = v$RDN_4516_out0 && v$_2746_out0;
assign v$G3_262_out0 = v$RDN_4517_out0 && v$_2747_out0;
assign v$G3_263_out0 = v$RDN_4518_out0 && v$_2748_out0;
assign v$G3_264_out0 = v$RDN_4519_out0 && v$_2749_out0;
assign v$G3_265_out0 = v$RDN_4520_out0 && v$_2750_out0;
assign v$G3_266_out0 = v$RDN_4521_out0 && v$_2751_out0;
assign v$G3_267_out0 = v$RDN_4522_out0 && v$_2752_out0;
assign v$G3_268_out0 = v$RDN_4523_out0 && v$_2753_out0;
assign v$G3_269_out0 = v$RDN_4524_out0 && v$_2754_out0;
assign v$G3_270_out0 = v$RDN_4525_out0 && v$_2755_out0;
assign v$G4_341_out0 = v$RDN_4496_out0 && v$_11098_out0;
assign v$G4_344_out0 = v$RDN_4499_out0 && v$_11101_out0;
assign v$G4_346_out0 = v$RDN_4501_out0 && v$_11103_out0;
assign v$G4_347_out0 = v$RDN_4502_out0 && v$_11104_out0;
assign v$G4_348_out0 = v$RDN_4503_out0 && v$_11105_out0;
assign v$G4_349_out0 = v$RDN_4504_out0 && v$_11106_out0;
assign v$G4_350_out0 = v$RDN_4505_out0 && v$_11107_out0;
assign v$G4_351_out0 = v$RDN_4506_out0 && v$_11108_out0;
assign v$G4_352_out0 = v$RDN_4507_out0 && v$_11109_out0;
assign v$G4_353_out0 = v$RDN_4508_out0 && v$_11110_out0;
assign v$G4_354_out0 = v$RDN_4509_out0 && v$_11111_out0;
assign v$G4_355_out0 = v$RDN_4510_out0 && v$_11112_out0;
assign v$G4_356_out0 = v$RDN_4511_out0 && v$_11113_out0;
assign v$G4_359_out0 = v$RDN_4514_out0 && v$_11116_out0;
assign v$G4_361_out0 = v$RDN_4516_out0 && v$_11118_out0;
assign v$G4_362_out0 = v$RDN_4517_out0 && v$_11119_out0;
assign v$G4_363_out0 = v$RDN_4518_out0 && v$_11120_out0;
assign v$G4_364_out0 = v$RDN_4519_out0 && v$_11121_out0;
assign v$G4_365_out0 = v$RDN_4520_out0 && v$_11122_out0;
assign v$G4_366_out0 = v$RDN_4521_out0 && v$_11123_out0;
assign v$G4_367_out0 = v$RDN_4522_out0 && v$_11124_out0;
assign v$G4_368_out0 = v$RDN_4523_out0 && v$_11125_out0;
assign v$G4_369_out0 = v$RDN_4524_out0 && v$_11126_out0;
assign v$G4_370_out0 = v$RDN_4525_out0 && v$_11127_out0;
assign v$_386_out0 = { v$G5_2783_out0,v$G6_8834_out0 };
assign v$_388_out0 = { v$G5_2785_out0,v$G6_8836_out0 };
assign v$_399_out0 = { v$G9_2895_out0,v$G10_2640_out0 };
assign v$_401_out0 = { v$G9_2897_out0,v$G10_2642_out0 };
assign v$G11_652_out0 = v$RD_13568_out0 && v$_3911_out0;
assign v$G11_653_out0 = v$RD_13569_out0 && v$_3912_out0;
assign v$G11_655_out0 = v$RD_13571_out0 && v$_3914_out0;
assign v$G11_667_out0 = v$RD_13583_out0 && v$_3926_out0;
assign v$G11_668_out0 = v$RD_13584_out0 && v$_3927_out0;
assign v$G11_670_out0 = v$RD_13586_out0 && v$_3929_out0;
assign v$2_1763_out0 = v$B_3946_out0[2:2];
assign v$2_1764_out0 = v$B_3947_out0[2:2];
assign v$G1_1909_out0 = v$RDN_4496_out0 && v$_568_out0;
assign v$G1_1912_out0 = v$RDN_4499_out0 && v$_571_out0;
assign v$G1_1914_out0 = v$RDN_4501_out0 && v$_573_out0;
assign v$G1_1915_out0 = v$RDN_4502_out0 && v$_574_out0;
assign v$G1_1916_out0 = v$RDN_4503_out0 && v$_575_out0;
assign v$G1_1917_out0 = v$RDN_4504_out0 && v$_576_out0;
assign v$G1_1918_out0 = v$RDN_4505_out0 && v$_577_out0;
assign v$G1_1919_out0 = v$RDN_4506_out0 && v$_578_out0;
assign v$G1_1920_out0 = v$RDN_4507_out0 && v$_579_out0;
assign v$G1_1921_out0 = v$RDN_4508_out0 && v$_580_out0;
assign v$G1_1922_out0 = v$RDN_4509_out0 && v$_581_out0;
assign v$G1_1923_out0 = v$RDN_4510_out0 && v$_582_out0;
assign v$G1_1924_out0 = v$RDN_4511_out0 && v$_583_out0;
assign v$G1_1927_out0 = v$RDN_4514_out0 && v$_586_out0;
assign v$G1_1929_out0 = v$RDN_4516_out0 && v$_588_out0;
assign v$G1_1930_out0 = v$RDN_4517_out0 && v$_589_out0;
assign v$G1_1931_out0 = v$RDN_4518_out0 && v$_590_out0;
assign v$G1_1932_out0 = v$RDN_4519_out0 && v$_591_out0;
assign v$G1_1933_out0 = v$RDN_4520_out0 && v$_592_out0;
assign v$G1_1934_out0 = v$RDN_4521_out0 && v$_593_out0;
assign v$G1_1935_out0 = v$RDN_4522_out0 && v$_594_out0;
assign v$G1_1936_out0 = v$RDN_4523_out0 && v$_595_out0;
assign v$G1_1937_out0 = v$RDN_4524_out0 && v$_596_out0;
assign v$G1_1938_out0 = v$RDN_4525_out0 && v$_597_out0;
assign v$G6_2116_out0 = v$RDN_4496_out0 && v$_13399_out0;
assign v$G6_2119_out0 = v$RDN_4499_out0 && v$_13402_out0;
assign v$G6_2121_out0 = v$RDN_4501_out0 && v$_13404_out0;
assign v$G6_2122_out0 = v$RDN_4502_out0 && v$_13405_out0;
assign v$G6_2123_out0 = v$RDN_4503_out0 && v$_13406_out0;
assign v$G6_2124_out0 = v$RDN_4504_out0 && v$_13407_out0;
assign v$G6_2125_out0 = v$RDN_4505_out0 && v$_13408_out0;
assign v$G6_2126_out0 = v$RDN_4506_out0 && v$_13409_out0;
assign v$G6_2127_out0 = v$RDN_4507_out0 && v$_13410_out0;
assign v$G6_2128_out0 = v$RDN_4508_out0 && v$_13411_out0;
assign v$G6_2129_out0 = v$RDN_4509_out0 && v$_13412_out0;
assign v$G6_2130_out0 = v$RDN_4510_out0 && v$_13413_out0;
assign v$G6_2131_out0 = v$RDN_4511_out0 && v$_13414_out0;
assign v$G6_2134_out0 = v$RDN_4514_out0 && v$_13417_out0;
assign v$G6_2136_out0 = v$RDN_4516_out0 && v$_13419_out0;
assign v$G6_2137_out0 = v$RDN_4517_out0 && v$_13420_out0;
assign v$G6_2138_out0 = v$RDN_4518_out0 && v$_13421_out0;
assign v$G6_2139_out0 = v$RDN_4519_out0 && v$_13422_out0;
assign v$G6_2140_out0 = v$RDN_4520_out0 && v$_13423_out0;
assign v$G6_2141_out0 = v$RDN_4521_out0 && v$_13424_out0;
assign v$G6_2142_out0 = v$RDN_4522_out0 && v$_13425_out0;
assign v$G6_2143_out0 = v$RDN_4523_out0 && v$_13426_out0;
assign v$G6_2144_out0 = v$RDN_4524_out0 && v$_13427_out0;
assign v$G6_2145_out0 = v$RDN_4525_out0 && v$_13428_out0;
assign v$G8_2472_out0 = v$RDN_4496_out0 && v$_2986_out0;
assign v$G8_2475_out0 = v$RDN_4499_out0 && v$_2989_out0;
assign v$G8_2477_out0 = v$RDN_4501_out0 && v$_2991_out0;
assign v$G8_2478_out0 = v$RDN_4502_out0 && v$_2992_out0;
assign v$G8_2479_out0 = v$RDN_4503_out0 && v$_2993_out0;
assign v$G8_2480_out0 = v$RDN_4504_out0 && v$_2994_out0;
assign v$G8_2481_out0 = v$RDN_4505_out0 && v$_2995_out0;
assign v$G8_2482_out0 = v$RDN_4506_out0 && v$_2996_out0;
assign v$G8_2483_out0 = v$RDN_4507_out0 && v$_2997_out0;
assign v$G8_2484_out0 = v$RDN_4508_out0 && v$_2998_out0;
assign v$G8_2485_out0 = v$RDN_4509_out0 && v$_2999_out0;
assign v$G8_2486_out0 = v$RDN_4510_out0 && v$_3000_out0;
assign v$G8_2487_out0 = v$RDN_4511_out0 && v$_3001_out0;
assign v$G8_2490_out0 = v$RDN_4514_out0 && v$_3004_out0;
assign v$G8_2492_out0 = v$RDN_4516_out0 && v$_3006_out0;
assign v$G8_2493_out0 = v$RDN_4517_out0 && v$_3007_out0;
assign v$G8_2494_out0 = v$RDN_4518_out0 && v$_3008_out0;
assign v$G8_2495_out0 = v$RDN_4519_out0 && v$_3009_out0;
assign v$G8_2496_out0 = v$RDN_4520_out0 && v$_3010_out0;
assign v$G8_2497_out0 = v$RDN_4521_out0 && v$_3011_out0;
assign v$G8_2498_out0 = v$RDN_4522_out0 && v$_3012_out0;
assign v$G8_2499_out0 = v$RDN_4523_out0 && v$_3013_out0;
assign v$G8_2500_out0 = v$RDN_4524_out0 && v$_3014_out0;
assign v$G8_2501_out0 = v$RDN_4525_out0 && v$_3015_out0;
assign v$_2649_out0 = { v$_2838_out0,v$G10_2632_out0 };
assign v$_2945_out0 = { v$G15_4654_out0,v$G16_10906_out0 };
assign v$_2947_out0 = { v$G15_4656_out0,v$G16_10908_out0 };
assign v$0_3022_out0 = v$B_3946_out0[0:0];
assign v$0_3023_out0 = v$B_3947_out0[0:0];
assign v$_3215_out0 = { v$G1_1879_out0,v$G2_1809_out0 };
assign v$_3217_out0 = { v$G1_1881_out0,v$G2_1811_out0 };
assign v$_3278_out0 = { v$G3_7087_out0,v$G4_2767_out0 };
assign v$_3280_out0 = { v$G3_7089_out0,v$G4_2769_out0 };
assign v$1_3817_out0 = v$B_3946_out0[1:1];
assign v$1_3818_out0 = v$B_3947_out0[1:1];
assign v$G2_4620_out0 = v$RDN_4496_out0 && v$_10874_out0;
assign v$G2_4623_out0 = v$RDN_4499_out0 && v$_10877_out0;
assign v$G2_4625_out0 = v$RDN_4501_out0 && v$_10879_out0;
assign v$G2_4626_out0 = v$RDN_4502_out0 && v$_10880_out0;
assign v$G2_4627_out0 = v$RDN_4503_out0 && v$_10881_out0;
assign v$G2_4628_out0 = v$RDN_4504_out0 && v$_10882_out0;
assign v$G2_4629_out0 = v$RDN_4505_out0 && v$_10883_out0;
assign v$G2_4630_out0 = v$RDN_4506_out0 && v$_10884_out0;
assign v$G2_4631_out0 = v$RDN_4507_out0 && v$_10885_out0;
assign v$G2_4632_out0 = v$RDN_4508_out0 && v$_10886_out0;
assign v$G2_4633_out0 = v$RDN_4509_out0 && v$_10887_out0;
assign v$G2_4634_out0 = v$RDN_4510_out0 && v$_10888_out0;
assign v$G2_4635_out0 = v$RDN_4511_out0 && v$_10889_out0;
assign v$G2_4638_out0 = v$RDN_4514_out0 && v$_10892_out0;
assign v$G2_4640_out0 = v$RDN_4516_out0 && v$_10894_out0;
assign v$G2_4641_out0 = v$RDN_4517_out0 && v$_10895_out0;
assign v$G2_4642_out0 = v$RDN_4518_out0 && v$_10896_out0;
assign v$G2_4643_out0 = v$RDN_4519_out0 && v$_10897_out0;
assign v$G2_4644_out0 = v$RDN_4520_out0 && v$_10898_out0;
assign v$G2_4645_out0 = v$RDN_4521_out0 && v$_10899_out0;
assign v$G2_4646_out0 = v$RDN_4522_out0 && v$_10900_out0;
assign v$G2_4647_out0 = v$RDN_4523_out0 && v$_10901_out0;
assign v$G2_4648_out0 = v$RDN_4524_out0 && v$_10902_out0;
assign v$G2_4649_out0 = v$RDN_4525_out0 && v$_10903_out0;
assign v$SIG$TO$SHIFT_5836_out0 = v$SIG$TO$SHIFT_10712_out0;
assign v$SIG$TO$SHIFT_5837_out0 = v$SIG$TO$SHIFT_10713_out0;
assign v$RD_5903_out0 = v$G16_13184_out0;
assign v$RD_5935_out0 = v$G16_13185_out0;
assign v$RD_5997_out0 = v$G16_13187_out0;
assign v$RD_6367_out0 = v$G16_13199_out0;
assign v$RD_6399_out0 = v$G16_13200_out0;
assign v$RD_6461_out0 = v$G16_13202_out0;
assign v$G10_6976_out0 = v$RD_13568_out0 && v$_2064_out0;
assign v$G10_6977_out0 = v$RD_13569_out0 && v$_2065_out0;
assign v$G10_6979_out0 = v$RD_13571_out0 && v$_2067_out0;
assign v$G10_6991_out0 = v$RD_13583_out0 && v$_2079_out0;
assign v$G10_6992_out0 = v$RD_13584_out0 && v$_2080_out0;
assign v$G10_6994_out0 = v$RD_13586_out0 && v$_2082_out0;
assign v$_7135_out0 = { v$G13_642_out0,v$G14_615_out0 };
assign v$_7137_out0 = { v$G13_644_out0,v$G14_617_out0 };
assign v$RD_7204_out0 = v$G5_10622_out0;
assign v$RD_7205_out0 = v$G2_4621_out0;
assign v$RD_7207_out0 = v$G9_10573_out0;
assign v$RD_7209_out0 = v$G1_1910_out0;
assign v$RD_7210_out0 = v$G4_342_out0;
assign v$RD_7211_out0 = v$G6_2117_out0;
assign v$RD_7212_out0 = v$G7_11263_out0;
assign v$RD_7214_out0 = v$G8_2473_out0;
assign v$RD_7215_out0 = v$G3_242_out0;
assign v$RD_7219_out0 = v$G5_10623_out0;
assign v$RD_7220_out0 = v$G2_4622_out0;
assign v$RD_7222_out0 = v$G9_10574_out0;
assign v$RD_7224_out0 = v$G1_1911_out0;
assign v$RD_7225_out0 = v$G4_343_out0;
assign v$RD_7226_out0 = v$G6_2118_out0;
assign v$RD_7227_out0 = v$G7_11264_out0;
assign v$RD_7229_out0 = v$G8_2474_out0;
assign v$RD_7230_out0 = v$G3_243_out0;
assign v$RD_7249_out0 = v$G5_10625_out0;
assign v$RD_7250_out0 = v$G2_4624_out0;
assign v$RD_7252_out0 = v$G9_10576_out0;
assign v$RD_7254_out0 = v$G1_1913_out0;
assign v$RD_7255_out0 = v$G4_345_out0;
assign v$RD_7256_out0 = v$G6_2120_out0;
assign v$RD_7257_out0 = v$G7_11266_out0;
assign v$RD_7259_out0 = v$G8_2476_out0;
assign v$RD_7260_out0 = v$G3_245_out0;
assign v$RD_7428_out0 = v$G5_10637_out0;
assign v$RD_7429_out0 = v$G2_4636_out0;
assign v$RD_7431_out0 = v$G9_10588_out0;
assign v$RD_7433_out0 = v$G1_1925_out0;
assign v$RD_7434_out0 = v$G4_357_out0;
assign v$RD_7435_out0 = v$G6_2132_out0;
assign v$RD_7436_out0 = v$G7_11278_out0;
assign v$RD_7438_out0 = v$G8_2488_out0;
assign v$RD_7439_out0 = v$G3_257_out0;
assign v$RD_7443_out0 = v$G5_10638_out0;
assign v$RD_7444_out0 = v$G2_4637_out0;
assign v$RD_7446_out0 = v$G9_10589_out0;
assign v$RD_7448_out0 = v$G1_1926_out0;
assign v$RD_7449_out0 = v$G4_358_out0;
assign v$RD_7450_out0 = v$G6_2133_out0;
assign v$RD_7451_out0 = v$G7_11279_out0;
assign v$RD_7453_out0 = v$G8_2489_out0;
assign v$RD_7454_out0 = v$G3_258_out0;
assign v$RD_7473_out0 = v$G5_10640_out0;
assign v$RD_7474_out0 = v$G2_4639_out0;
assign v$RD_7476_out0 = v$G9_10591_out0;
assign v$RD_7478_out0 = v$G1_1928_out0;
assign v$RD_7479_out0 = v$G4_360_out0;
assign v$RD_7480_out0 = v$G6_2135_out0;
assign v$RD_7481_out0 = v$G7_11281_out0;
assign v$RD_7483_out0 = v$G8_2491_out0;
assign v$RD_7484_out0 = v$G3_260_out0;
assign v$SUBNORMAL_8808_out0 = v$EQ1_6956_out0;
assign v$SUBNORMAL_8809_out0 = v$EQ1_6957_out0;
assign v$IN_10403_out0 = v$OUT_1136_out0;
assign v$IN_10404_out0 = v$OUT_1137_out0;
assign v$_10456_out0 = { v$_174_out0,v$G15_1815_out0 };
assign v$_10458_out0 = { v$_176_out0,v$G15_1817_out0 };
assign v$G9_10572_out0 = v$RDN_4496_out0 && v$_3961_out0;
assign v$G9_10575_out0 = v$RDN_4499_out0 && v$_3964_out0;
assign v$G9_10577_out0 = v$RDN_4501_out0 && v$_3966_out0;
assign v$G9_10578_out0 = v$RDN_4502_out0 && v$_3967_out0;
assign v$G9_10579_out0 = v$RDN_4503_out0 && v$_3968_out0;
assign v$G9_10580_out0 = v$RDN_4504_out0 && v$_3969_out0;
assign v$G9_10581_out0 = v$RDN_4505_out0 && v$_3970_out0;
assign v$G9_10582_out0 = v$RDN_4506_out0 && v$_3971_out0;
assign v$G9_10583_out0 = v$RDN_4507_out0 && v$_3972_out0;
assign v$G9_10584_out0 = v$RDN_4508_out0 && v$_3973_out0;
assign v$G9_10585_out0 = v$RDN_4509_out0 && v$_3974_out0;
assign v$G9_10586_out0 = v$RDN_4510_out0 && v$_3975_out0;
assign v$G9_10587_out0 = v$RDN_4511_out0 && v$_3976_out0;
assign v$G9_10590_out0 = v$RDN_4514_out0 && v$_3979_out0;
assign v$G9_10592_out0 = v$RDN_4516_out0 && v$_3981_out0;
assign v$G9_10593_out0 = v$RDN_4517_out0 && v$_3982_out0;
assign v$G9_10594_out0 = v$RDN_4518_out0 && v$_3983_out0;
assign v$G9_10595_out0 = v$RDN_4519_out0 && v$_3984_out0;
assign v$G9_10596_out0 = v$RDN_4520_out0 && v$_3985_out0;
assign v$G9_10597_out0 = v$RDN_4521_out0 && v$_3986_out0;
assign v$G9_10598_out0 = v$RDN_4522_out0 && v$_3987_out0;
assign v$G9_10599_out0 = v$RDN_4523_out0 && v$_3988_out0;
assign v$G9_10600_out0 = v$RDN_4524_out0 && v$_3989_out0;
assign v$G9_10601_out0 = v$RDN_4525_out0 && v$_3990_out0;
assign v$G5_10621_out0 = v$RDN_4496_out0 && v$_503_out0;
assign v$G5_10624_out0 = v$RDN_4499_out0 && v$_506_out0;
assign v$G5_10626_out0 = v$RDN_4501_out0 && v$_508_out0;
assign v$G5_10627_out0 = v$RDN_4502_out0 && v$_509_out0;
assign v$G5_10628_out0 = v$RDN_4503_out0 && v$_510_out0;
assign v$G5_10629_out0 = v$RDN_4504_out0 && v$_511_out0;
assign v$G5_10630_out0 = v$RDN_4505_out0 && v$_512_out0;
assign v$G5_10631_out0 = v$RDN_4506_out0 && v$_513_out0;
assign v$G5_10632_out0 = v$RDN_4507_out0 && v$_514_out0;
assign v$G5_10633_out0 = v$RDN_4508_out0 && v$_515_out0;
assign v$G5_10634_out0 = v$RDN_4509_out0 && v$_516_out0;
assign v$G5_10635_out0 = v$RDN_4510_out0 && v$_517_out0;
assign v$G5_10636_out0 = v$RDN_4511_out0 && v$_518_out0;
assign v$G5_10639_out0 = v$RDN_4514_out0 && v$_521_out0;
assign v$G5_10641_out0 = v$RDN_4516_out0 && v$_523_out0;
assign v$G5_10642_out0 = v$RDN_4517_out0 && v$_524_out0;
assign v$G5_10643_out0 = v$RDN_4518_out0 && v$_525_out0;
assign v$G5_10644_out0 = v$RDN_4519_out0 && v$_526_out0;
assign v$G5_10645_out0 = v$RDN_4520_out0 && v$_527_out0;
assign v$G5_10646_out0 = v$RDN_4521_out0 && v$_528_out0;
assign v$G5_10647_out0 = v$RDN_4522_out0 && v$_529_out0;
assign v$G5_10648_out0 = v$RDN_4523_out0 && v$_530_out0;
assign v$G5_10649_out0 = v$RDN_4524_out0 && v$_531_out0;
assign v$G5_10650_out0 = v$RDN_4525_out0 && v$_532_out0;
assign v$G7_11262_out0 = v$RDN_4496_out0 && v$_10409_out0;
assign v$G7_11265_out0 = v$RDN_4499_out0 && v$_10412_out0;
assign v$G7_11267_out0 = v$RDN_4501_out0 && v$_10414_out0;
assign v$G7_11268_out0 = v$RDN_4502_out0 && v$_10415_out0;
assign v$G7_11269_out0 = v$RDN_4503_out0 && v$_10416_out0;
assign v$G7_11270_out0 = v$RDN_4504_out0 && v$_10417_out0;
assign v$G7_11271_out0 = v$RDN_4505_out0 && v$_10418_out0;
assign v$G7_11272_out0 = v$RDN_4506_out0 && v$_10419_out0;
assign v$G7_11273_out0 = v$RDN_4507_out0 && v$_10420_out0;
assign v$G7_11274_out0 = v$RDN_4508_out0 && v$_10421_out0;
assign v$G7_11275_out0 = v$RDN_4509_out0 && v$_10422_out0;
assign v$G7_11276_out0 = v$RDN_4510_out0 && v$_10423_out0;
assign v$G7_11277_out0 = v$RDN_4511_out0 && v$_10424_out0;
assign v$G7_11280_out0 = v$RDN_4514_out0 && v$_10427_out0;
assign v$G7_11282_out0 = v$RDN_4516_out0 && v$_10429_out0;
assign v$G7_11283_out0 = v$RDN_4517_out0 && v$_10430_out0;
assign v$G7_11284_out0 = v$RDN_4518_out0 && v$_10431_out0;
assign v$G7_11285_out0 = v$RDN_4519_out0 && v$_10432_out0;
assign v$G7_11286_out0 = v$RDN_4520_out0 && v$_10433_out0;
assign v$G7_11287_out0 = v$RDN_4521_out0 && v$_10434_out0;
assign v$G7_11288_out0 = v$RDN_4522_out0 && v$_10435_out0;
assign v$G7_11289_out0 = v$RDN_4523_out0 && v$_10436_out0;
assign v$G7_11290_out0 = v$RDN_4524_out0 && v$_10437_out0;
assign v$G7_11291_out0 = v$RDN_4525_out0 && v$_10438_out0;
assign v$G16_13183_out0 = v$RDN_4496_out0 && v$_11001_out0;
assign v$G16_13186_out0 = v$RDN_4499_out0 && v$_11004_out0;
assign v$G16_13188_out0 = v$RDN_4501_out0 && v$_11006_out0;
assign v$G16_13189_out0 = v$RDN_4502_out0 && v$_11007_out0;
assign v$G16_13190_out0 = v$RDN_4503_out0 && v$_11008_out0;
assign v$G16_13191_out0 = v$RDN_4504_out0 && v$_11009_out0;
assign v$G16_13192_out0 = v$RDN_4505_out0 && v$_11010_out0;
assign v$G16_13193_out0 = v$RDN_4506_out0 && v$_11011_out0;
assign v$G16_13194_out0 = v$RDN_4507_out0 && v$_11012_out0;
assign v$G16_13195_out0 = v$RDN_4508_out0 && v$_11013_out0;
assign v$G16_13196_out0 = v$RDN_4509_out0 && v$_11014_out0;
assign v$G16_13197_out0 = v$RDN_4510_out0 && v$_11015_out0;
assign v$G16_13198_out0 = v$RDN_4511_out0 && v$_11016_out0;
assign v$G16_13201_out0 = v$RDN_4514_out0 && v$_11019_out0;
assign v$G16_13203_out0 = v$RDN_4516_out0 && v$_11021_out0;
assign v$G16_13204_out0 = v$RDN_4517_out0 && v$_11022_out0;
assign v$G16_13205_out0 = v$RDN_4518_out0 && v$_11023_out0;
assign v$G16_13206_out0 = v$RDN_4519_out0 && v$_11024_out0;
assign v$G16_13207_out0 = v$RDN_4520_out0 && v$_11025_out0;
assign v$G16_13208_out0 = v$RDN_4521_out0 && v$_11026_out0;
assign v$G16_13209_out0 = v$RDN_4522_out0 && v$_11027_out0;
assign v$G16_13210_out0 = v$RDN_4523_out0 && v$_11028_out0;
assign v$G16_13211_out0 = v$RDN_4524_out0 && v$_11029_out0;
assign v$G16_13212_out0 = v$RDN_4525_out0 && v$_11030_out0;
assign v$G12_13222_out0 = v$RD_13568_out0 && v$_2274_out0;
assign v$G12_13223_out0 = v$RD_13569_out0 && v$_2275_out0;
assign v$G12_13225_out0 = v$RD_13571_out0 && v$_2277_out0;
assign v$G12_13237_out0 = v$RD_13583_out0 && v$_2289_out0;
assign v$G12_13238_out0 = v$RD_13584_out0 && v$_2290_out0;
assign v$G12_13240_out0 = v$RD_13586_out0 && v$_2292_out0;
assign v$_13261_out0 = { v$G11_2937_out0,v$G12_10688_out0 };
assign v$_13263_out0 = { v$G11_2939_out0,v$G12_10690_out0 };
assign v$G13_13353_out0 = v$RD_13568_out0 && v$_13716_out0;
assign v$G13_13354_out0 = v$RD_13569_out0 && v$_13717_out0;
assign v$G13_13356_out0 = v$RD_13571_out0 && v$_13719_out0;
assign v$G13_13368_out0 = v$RD_13583_out0 && v$_13731_out0;
assign v$G13_13369_out0 = v$RD_13584_out0 && v$_13732_out0;
assign v$G13_13371_out0 = v$RD_13586_out0 && v$_13734_out0;
assign v$EXP1_13488_out0 = v$EQ2_11254_out0;
assign v$EXP1_13489_out0 = v$EQ2_11255_out0;
assign v$RD_13567_out0 = v$RDN_4496_out0;
assign v$RD_13570_out0 = v$RDN_4499_out0;
assign v$RD_13572_out0 = v$RDN_4501_out0;
assign v$RD_13573_out0 = v$RDN_4502_out0;
assign v$RD_13574_out0 = v$RDN_4503_out0;
assign v$RD_13575_out0 = v$RDN_4504_out0;
assign v$RD_13576_out0 = v$RDN_4505_out0;
assign v$RD_13577_out0 = v$RDN_4506_out0;
assign v$RD_13578_out0 = v$RDN_4507_out0;
assign v$RD_13579_out0 = v$RDN_4508_out0;
assign v$RD_13580_out0 = v$RDN_4509_out0;
assign v$RD_13581_out0 = v$RDN_4510_out0;
assign v$RD_13582_out0 = v$RDN_4511_out0;
assign v$RD_13585_out0 = v$RDN_4514_out0;
assign v$RD_13587_out0 = v$RDN_4516_out0;
assign v$RD_13588_out0 = v$RDN_4517_out0;
assign v$RD_13589_out0 = v$RDN_4518_out0;
assign v$RD_13590_out0 = v$RDN_4519_out0;
assign v$RD_13591_out0 = v$RDN_4520_out0;
assign v$RD_13592_out0 = v$RDN_4521_out0;
assign v$RD_13593_out0 = v$RDN_4522_out0;
assign v$RD_13594_out0 = v$RDN_4523_out0;
assign v$RD_13595_out0 = v$RDN_4524_out0;
assign v$RD_13596_out0 = v$RDN_4525_out0;
assign v$3_13619_out0 = v$B_3946_out0[3:3];
assign v$3_13620_out0 = v$B_3947_out0[3:3];
assign v$G14_13673_out0 = v$RD_13568_out0 && v$_6831_out0;
assign v$G14_13674_out0 = v$RD_13569_out0 && v$_6832_out0;
assign v$G14_13676_out0 = v$RD_13571_out0 && v$_6834_out0;
assign v$G14_13688_out0 = v$RD_13583_out0 && v$_6846_out0;
assign v$G14_13689_out0 = v$RD_13584_out0 && v$_6847_out0;
assign v$G14_13691_out0 = v$RD_13586_out0 && v$_6849_out0;
assign v$_13770_out0 = { v$G7_8655_out0,v$G8_548_out0 };
assign v$_13772_out0 = { v$G7_8657_out0,v$G8_550_out0 };
assign v$_113_out0 = { v$_386_out0,v$_13770_out0 };
assign v$_115_out0 = { v$_388_out0,v$_13772_out0 };
assign v$G15_132_out0 = v$RD_13567_out0 && v$_1975_out0;
assign v$G15_135_out0 = v$RD_13570_out0 && v$_1978_out0;
assign v$G15_137_out0 = v$RD_13572_out0 && v$_1980_out0;
assign v$G15_138_out0 = v$RD_13573_out0 && v$_1981_out0;
assign v$G15_139_out0 = v$RD_13574_out0 && v$_1982_out0;
assign v$G15_140_out0 = v$RD_13575_out0 && v$_1983_out0;
assign v$G15_141_out0 = v$RD_13576_out0 && v$_1984_out0;
assign v$G15_142_out0 = v$RD_13577_out0 && v$_1985_out0;
assign v$G15_143_out0 = v$RD_13578_out0 && v$_1986_out0;
assign v$G15_144_out0 = v$RD_13579_out0 && v$_1987_out0;
assign v$G15_145_out0 = v$RD_13580_out0 && v$_1988_out0;
assign v$G15_146_out0 = v$RD_13581_out0 && v$_1989_out0;
assign v$G15_147_out0 = v$RD_13582_out0 && v$_1990_out0;
assign v$G15_150_out0 = v$RD_13585_out0 && v$_1993_out0;
assign v$G15_152_out0 = v$RD_13587_out0 && v$_1995_out0;
assign v$G15_153_out0 = v$RD_13588_out0 && v$_1996_out0;
assign v$G15_154_out0 = v$RD_13589_out0 && v$_1997_out0;
assign v$G15_155_out0 = v$RD_13590_out0 && v$_1998_out0;
assign v$G15_156_out0 = v$RD_13591_out0 && v$_1999_out0;
assign v$G15_157_out0 = v$RD_13592_out0 && v$_2000_out0;
assign v$G15_158_out0 = v$RD_13593_out0 && v$_2001_out0;
assign v$G15_159_out0 = v$RD_13594_out0 && v$_2002_out0;
assign v$G15_160_out0 = v$RD_13595_out0 && v$_2003_out0;
assign v$G15_161_out0 = v$RD_13596_out0 && v$_2004_out0;
assign v$_449_out0 = { v$_7135_out0,v$_2945_out0 };
assign v$_451_out0 = { v$_7137_out0,v$_2947_out0 };
assign v$G5_638_out0 = ! v$EXP1_13488_out0;
assign v$G5_639_out0 = ! v$EXP1_13489_out0;
assign v$G11_651_out0 = v$RD_13567_out0 && v$_3910_out0;
assign v$G11_654_out0 = v$RD_13570_out0 && v$_3913_out0;
assign v$G11_656_out0 = v$RD_13572_out0 && v$_3915_out0;
assign v$G11_657_out0 = v$RD_13573_out0 && v$_3916_out0;
assign v$G11_658_out0 = v$RD_13574_out0 && v$_3917_out0;
assign v$G11_659_out0 = v$RD_13575_out0 && v$_3918_out0;
assign v$G11_660_out0 = v$RD_13576_out0 && v$_3919_out0;
assign v$G11_661_out0 = v$RD_13577_out0 && v$_3920_out0;
assign v$G11_662_out0 = v$RD_13578_out0 && v$_3921_out0;
assign v$G11_663_out0 = v$RD_13579_out0 && v$_3922_out0;
assign v$G11_664_out0 = v$RD_13580_out0 && v$_3923_out0;
assign v$G11_665_out0 = v$RD_13581_out0 && v$_3924_out0;
assign v$G11_666_out0 = v$RD_13582_out0 && v$_3925_out0;
assign v$G11_669_out0 = v$RD_13585_out0 && v$_3928_out0;
assign v$G11_671_out0 = v$RD_13587_out0 && v$_3930_out0;
assign v$G11_672_out0 = v$RD_13588_out0 && v$_3931_out0;
assign v$G11_673_out0 = v$RD_13589_out0 && v$_3932_out0;
assign v$G11_674_out0 = v$RD_13590_out0 && v$_3933_out0;
assign v$G11_675_out0 = v$RD_13591_out0 && v$_3934_out0;
assign v$G11_676_out0 = v$RD_13592_out0 && v$_3935_out0;
assign v$G11_677_out0 = v$RD_13593_out0 && v$_3936_out0;
assign v$G11_678_out0 = v$RD_13594_out0 && v$_3937_out0;
assign v$G11_679_out0 = v$RD_13595_out0 && v$_3938_out0;
assign v$G11_680_out0 = v$RD_13596_out0 && v$_3939_out0;
assign v$_1212_out0 = { v$_10456_out0,v$G16_11035_out0 };
assign v$_1214_out0 = { v$_10458_out0,v$G16_11037_out0 };
assign v$_2345_out0 = { v$_399_out0,v$_13261_out0 };
assign v$_2347_out0 = { v$_401_out0,v$_13263_out0 };
assign v$_4733_out0 = { v$_2649_out0,v$G11_2550_out0 };
assign v$RD_5874_out0 = v$G16_13183_out0;
assign v$RD_5897_out0 = v$RD_7204_out0;
assign v$RD_5899_out0 = v$RD_7205_out0;
assign v$RD_5904_out0 = v$G15_133_out0;
assign v$RD_5905_out0 = v$RD_7207_out0;
assign v$RD_5909_out0 = v$RD_7209_out0;
assign v$RD_5911_out0 = v$RD_7210_out0;
assign v$RD_5913_out0 = v$RD_7211_out0;
assign v$RD_5915_out0 = v$RD_7212_out0;
assign v$RD_5919_out0 = v$RD_7214_out0;
assign v$RD_5921_out0 = v$RD_7215_out0;
assign v$RD_5929_out0 = v$RD_7219_out0;
assign v$RD_5931_out0 = v$RD_7220_out0;
assign v$RD_5936_out0 = v$RD_7222_out0;
assign v$RD_5940_out0 = v$RD_7224_out0;
assign v$RD_5942_out0 = v$RD_7225_out0;
assign v$RD_5944_out0 = v$RD_7226_out0;
assign v$RD_5946_out0 = v$RD_7227_out0;
assign v$RD_5950_out0 = v$RD_7229_out0;
assign v$RD_5952_out0 = v$RD_7230_out0;
assign v$RD_5966_out0 = v$G16_13186_out0;
assign v$RD_5991_out0 = v$RD_7249_out0;
assign v$RD_5993_out0 = v$RD_7250_out0;
assign v$RD_5998_out0 = v$RD_7252_out0;
assign v$RD_6002_out0 = v$RD_7254_out0;
assign v$RD_6004_out0 = v$RD_7255_out0;
assign v$RD_6006_out0 = v$RD_7256_out0;
assign v$RD_6008_out0 = v$RD_7257_out0;
assign v$RD_6012_out0 = v$RD_7259_out0;
assign v$RD_6014_out0 = v$RD_7260_out0;
assign v$RD_6028_out0 = v$G16_13188_out0;
assign v$RD_6059_out0 = v$G16_13189_out0;
assign v$RD_6090_out0 = v$G16_13190_out0;
assign v$RD_6121_out0 = v$G16_13191_out0;
assign v$RD_6152_out0 = v$G16_13192_out0;
assign v$RD_6183_out0 = v$G16_13193_out0;
assign v$RD_6214_out0 = v$G16_13194_out0;
assign v$RD_6245_out0 = v$G16_13195_out0;
assign v$RD_6276_out0 = v$G16_13196_out0;
assign v$RD_6307_out0 = v$G16_13197_out0;
assign v$RD_6338_out0 = v$G16_13198_out0;
assign v$RD_6361_out0 = v$RD_7428_out0;
assign v$RD_6363_out0 = v$RD_7429_out0;
assign v$RD_6368_out0 = v$G15_148_out0;
assign v$RD_6369_out0 = v$RD_7431_out0;
assign v$RD_6373_out0 = v$RD_7433_out0;
assign v$RD_6375_out0 = v$RD_7434_out0;
assign v$RD_6377_out0 = v$RD_7435_out0;
assign v$RD_6379_out0 = v$RD_7436_out0;
assign v$RD_6383_out0 = v$RD_7438_out0;
assign v$RD_6385_out0 = v$RD_7439_out0;
assign v$RD_6393_out0 = v$RD_7443_out0;
assign v$RD_6395_out0 = v$RD_7444_out0;
assign v$RD_6400_out0 = v$RD_7446_out0;
assign v$RD_6404_out0 = v$RD_7448_out0;
assign v$RD_6406_out0 = v$RD_7449_out0;
assign v$RD_6408_out0 = v$RD_7450_out0;
assign v$RD_6410_out0 = v$RD_7451_out0;
assign v$RD_6414_out0 = v$RD_7453_out0;
assign v$RD_6416_out0 = v$RD_7454_out0;
assign v$RD_6430_out0 = v$G16_13201_out0;
assign v$RD_6455_out0 = v$RD_7473_out0;
assign v$RD_6457_out0 = v$RD_7474_out0;
assign v$RD_6462_out0 = v$RD_7476_out0;
assign v$RD_6466_out0 = v$RD_7478_out0;
assign v$RD_6468_out0 = v$RD_7479_out0;
assign v$RD_6470_out0 = v$RD_7480_out0;
assign v$RD_6472_out0 = v$RD_7481_out0;
assign v$RD_6476_out0 = v$RD_7483_out0;
assign v$RD_6478_out0 = v$RD_7484_out0;
assign v$RD_6492_out0 = v$G16_13203_out0;
assign v$RD_6523_out0 = v$G16_13204_out0;
assign v$RD_6554_out0 = v$G16_13205_out0;
assign v$RD_6585_out0 = v$G16_13206_out0;
assign v$RD_6616_out0 = v$G16_13207_out0;
assign v$RD_6647_out0 = v$G16_13208_out0;
assign v$RD_6678_out0 = v$G16_13209_out0;
assign v$RD_6709_out0 = v$G16_13210_out0;
assign v$RD_6740_out0 = v$G16_13211_out0;
assign v$RD_6771_out0 = v$G16_13212_out0;
assign v$G10_6975_out0 = v$RD_13567_out0 && v$_2063_out0;
assign v$G10_6978_out0 = v$RD_13570_out0 && v$_2066_out0;
assign v$G10_6980_out0 = v$RD_13572_out0 && v$_2068_out0;
assign v$G10_6981_out0 = v$RD_13573_out0 && v$_2069_out0;
assign v$G10_6982_out0 = v$RD_13574_out0 && v$_2070_out0;
assign v$G10_6983_out0 = v$RD_13575_out0 && v$_2071_out0;
assign v$G10_6984_out0 = v$RD_13576_out0 && v$_2072_out0;
assign v$G10_6985_out0 = v$RD_13577_out0 && v$_2073_out0;
assign v$G10_6986_out0 = v$RD_13578_out0 && v$_2074_out0;
assign v$G10_6987_out0 = v$RD_13579_out0 && v$_2075_out0;
assign v$G10_6988_out0 = v$RD_13580_out0 && v$_2076_out0;
assign v$G10_6989_out0 = v$RD_13581_out0 && v$_2077_out0;
assign v$G10_6990_out0 = v$RD_13582_out0 && v$_2078_out0;
assign v$G10_6993_out0 = v$RD_13585_out0 && v$_2081_out0;
assign v$G10_6995_out0 = v$RD_13587_out0 && v$_2083_out0;
assign v$G10_6996_out0 = v$RD_13588_out0 && v$_2084_out0;
assign v$G10_6997_out0 = v$RD_13589_out0 && v$_2085_out0;
assign v$G10_6998_out0 = v$RD_13590_out0 && v$_2086_out0;
assign v$G10_6999_out0 = v$RD_13591_out0 && v$_2087_out0;
assign v$G10_7000_out0 = v$RD_13592_out0 && v$_2088_out0;
assign v$G10_7001_out0 = v$RD_13593_out0 && v$_2089_out0;
assign v$G10_7002_out0 = v$RD_13594_out0 && v$_2090_out0;
assign v$G10_7003_out0 = v$RD_13595_out0 && v$_2091_out0;
assign v$G10_7004_out0 = v$RD_13596_out0 && v$_2092_out0;
assign v$RD_7190_out0 = v$G5_10621_out0;
assign v$RD_7191_out0 = v$G2_4620_out0;
assign v$RD_7193_out0 = v$G9_10572_out0;
assign v$RD_7195_out0 = v$G1_1909_out0;
assign v$RD_7196_out0 = v$G4_341_out0;
assign v$RD_7197_out0 = v$G6_2116_out0;
assign v$RD_7198_out0 = v$G7_11262_out0;
assign v$RD_7200_out0 = v$G8_2472_out0;
assign v$RD_7201_out0 = v$G3_241_out0;
assign v$RD_7202_out0 = v$G12_13222_out0;
assign v$RD_7203_out0 = v$G14_13673_out0;
assign v$RD_7206_out0 = v$G13_13353_out0;
assign v$RD_7208_out0 = v$G10_6976_out0;
assign v$RD_7213_out0 = v$G11_652_out0;
assign v$RD_7216_out0 = v$G12_13223_out0;
assign v$RD_7217_out0 = v$G14_13674_out0;
assign v$RD_7218_out0 = v$G15_134_out0;
assign v$RD_7221_out0 = v$G13_13354_out0;
assign v$RD_7223_out0 = v$G10_6977_out0;
assign v$RD_7228_out0 = v$G11_653_out0;
assign v$RD_7234_out0 = v$G5_10624_out0;
assign v$RD_7235_out0 = v$G2_4623_out0;
assign v$RD_7237_out0 = v$G9_10575_out0;
assign v$RD_7239_out0 = v$G1_1912_out0;
assign v$RD_7240_out0 = v$G4_344_out0;
assign v$RD_7241_out0 = v$G6_2119_out0;
assign v$RD_7242_out0 = v$G7_11265_out0;
assign v$RD_7244_out0 = v$G8_2475_out0;
assign v$RD_7245_out0 = v$G3_244_out0;
assign v$RD_7246_out0 = v$G12_13225_out0;
assign v$RD_7247_out0 = v$G14_13676_out0;
assign v$RD_7248_out0 = v$G15_136_out0;
assign v$RD_7251_out0 = v$G13_13356_out0;
assign v$RD_7253_out0 = v$G10_6979_out0;
assign v$RD_7258_out0 = v$G11_655_out0;
assign v$RD_7264_out0 = v$G5_10626_out0;
assign v$RD_7265_out0 = v$G2_4625_out0;
assign v$RD_7267_out0 = v$G9_10577_out0;
assign v$RD_7269_out0 = v$G1_1914_out0;
assign v$RD_7270_out0 = v$G4_346_out0;
assign v$RD_7271_out0 = v$G6_2121_out0;
assign v$RD_7272_out0 = v$G7_11267_out0;
assign v$RD_7274_out0 = v$G8_2477_out0;
assign v$RD_7275_out0 = v$G3_246_out0;
assign v$RD_7279_out0 = v$G5_10627_out0;
assign v$RD_7280_out0 = v$G2_4626_out0;
assign v$RD_7282_out0 = v$G9_10578_out0;
assign v$RD_7284_out0 = v$G1_1915_out0;
assign v$RD_7285_out0 = v$G4_347_out0;
assign v$RD_7286_out0 = v$G6_2122_out0;
assign v$RD_7287_out0 = v$G7_11268_out0;
assign v$RD_7289_out0 = v$G8_2478_out0;
assign v$RD_7290_out0 = v$G3_247_out0;
assign v$RD_7294_out0 = v$G5_10628_out0;
assign v$RD_7295_out0 = v$G2_4627_out0;
assign v$RD_7297_out0 = v$G9_10579_out0;
assign v$RD_7299_out0 = v$G1_1916_out0;
assign v$RD_7300_out0 = v$G4_348_out0;
assign v$RD_7301_out0 = v$G6_2123_out0;
assign v$RD_7302_out0 = v$G7_11269_out0;
assign v$RD_7304_out0 = v$G8_2479_out0;
assign v$RD_7305_out0 = v$G3_248_out0;
assign v$RD_7309_out0 = v$G5_10629_out0;
assign v$RD_7310_out0 = v$G2_4628_out0;
assign v$RD_7312_out0 = v$G9_10580_out0;
assign v$RD_7314_out0 = v$G1_1917_out0;
assign v$RD_7315_out0 = v$G4_349_out0;
assign v$RD_7316_out0 = v$G6_2124_out0;
assign v$RD_7317_out0 = v$G7_11270_out0;
assign v$RD_7319_out0 = v$G8_2480_out0;
assign v$RD_7320_out0 = v$G3_249_out0;
assign v$RD_7324_out0 = v$G5_10630_out0;
assign v$RD_7325_out0 = v$G2_4629_out0;
assign v$RD_7327_out0 = v$G9_10581_out0;
assign v$RD_7329_out0 = v$G1_1918_out0;
assign v$RD_7330_out0 = v$G4_350_out0;
assign v$RD_7331_out0 = v$G6_2125_out0;
assign v$RD_7332_out0 = v$G7_11271_out0;
assign v$RD_7334_out0 = v$G8_2481_out0;
assign v$RD_7335_out0 = v$G3_250_out0;
assign v$RD_7339_out0 = v$G5_10631_out0;
assign v$RD_7340_out0 = v$G2_4630_out0;
assign v$RD_7342_out0 = v$G9_10582_out0;
assign v$RD_7344_out0 = v$G1_1919_out0;
assign v$RD_7345_out0 = v$G4_351_out0;
assign v$RD_7346_out0 = v$G6_2126_out0;
assign v$RD_7347_out0 = v$G7_11272_out0;
assign v$RD_7349_out0 = v$G8_2482_out0;
assign v$RD_7350_out0 = v$G3_251_out0;
assign v$RD_7354_out0 = v$G5_10632_out0;
assign v$RD_7355_out0 = v$G2_4631_out0;
assign v$RD_7357_out0 = v$G9_10583_out0;
assign v$RD_7359_out0 = v$G1_1920_out0;
assign v$RD_7360_out0 = v$G4_352_out0;
assign v$RD_7361_out0 = v$G6_2127_out0;
assign v$RD_7362_out0 = v$G7_11273_out0;
assign v$RD_7364_out0 = v$G8_2483_out0;
assign v$RD_7365_out0 = v$G3_252_out0;
assign v$RD_7369_out0 = v$G5_10633_out0;
assign v$RD_7370_out0 = v$G2_4632_out0;
assign v$RD_7372_out0 = v$G9_10584_out0;
assign v$RD_7374_out0 = v$G1_1921_out0;
assign v$RD_7375_out0 = v$G4_353_out0;
assign v$RD_7376_out0 = v$G6_2128_out0;
assign v$RD_7377_out0 = v$G7_11274_out0;
assign v$RD_7379_out0 = v$G8_2484_out0;
assign v$RD_7380_out0 = v$G3_253_out0;
assign v$RD_7384_out0 = v$G5_10634_out0;
assign v$RD_7385_out0 = v$G2_4633_out0;
assign v$RD_7387_out0 = v$G9_10585_out0;
assign v$RD_7389_out0 = v$G1_1922_out0;
assign v$RD_7390_out0 = v$G4_354_out0;
assign v$RD_7391_out0 = v$G6_2129_out0;
assign v$RD_7392_out0 = v$G7_11275_out0;
assign v$RD_7394_out0 = v$G8_2485_out0;
assign v$RD_7395_out0 = v$G3_254_out0;
assign v$RD_7399_out0 = v$G5_10635_out0;
assign v$RD_7400_out0 = v$G2_4634_out0;
assign v$RD_7402_out0 = v$G9_10586_out0;
assign v$RD_7404_out0 = v$G1_1923_out0;
assign v$RD_7405_out0 = v$G4_355_out0;
assign v$RD_7406_out0 = v$G6_2130_out0;
assign v$RD_7407_out0 = v$G7_11276_out0;
assign v$RD_7409_out0 = v$G8_2486_out0;
assign v$RD_7410_out0 = v$G3_255_out0;
assign v$RD_7414_out0 = v$G5_10636_out0;
assign v$RD_7415_out0 = v$G2_4635_out0;
assign v$RD_7417_out0 = v$G9_10587_out0;
assign v$RD_7419_out0 = v$G1_1924_out0;
assign v$RD_7420_out0 = v$G4_356_out0;
assign v$RD_7421_out0 = v$G6_2131_out0;
assign v$RD_7422_out0 = v$G7_11277_out0;
assign v$RD_7424_out0 = v$G8_2487_out0;
assign v$RD_7425_out0 = v$G3_256_out0;
assign v$RD_7426_out0 = v$G12_13237_out0;
assign v$RD_7427_out0 = v$G14_13688_out0;
assign v$RD_7430_out0 = v$G13_13368_out0;
assign v$RD_7432_out0 = v$G10_6991_out0;
assign v$RD_7437_out0 = v$G11_667_out0;
assign v$RD_7440_out0 = v$G12_13238_out0;
assign v$RD_7441_out0 = v$G14_13689_out0;
assign v$RD_7442_out0 = v$G15_149_out0;
assign v$RD_7445_out0 = v$G13_13369_out0;
assign v$RD_7447_out0 = v$G10_6992_out0;
assign v$RD_7452_out0 = v$G11_668_out0;
assign v$RD_7458_out0 = v$G5_10639_out0;
assign v$RD_7459_out0 = v$G2_4638_out0;
assign v$RD_7461_out0 = v$G9_10590_out0;
assign v$RD_7463_out0 = v$G1_1927_out0;
assign v$RD_7464_out0 = v$G4_359_out0;
assign v$RD_7465_out0 = v$G6_2134_out0;
assign v$RD_7466_out0 = v$G7_11280_out0;
assign v$RD_7468_out0 = v$G8_2490_out0;
assign v$RD_7469_out0 = v$G3_259_out0;
assign v$RD_7470_out0 = v$G12_13240_out0;
assign v$RD_7471_out0 = v$G14_13691_out0;
assign v$RD_7472_out0 = v$G15_151_out0;
assign v$RD_7475_out0 = v$G13_13371_out0;
assign v$RD_7477_out0 = v$G10_6994_out0;
assign v$RD_7482_out0 = v$G11_670_out0;
assign v$RD_7488_out0 = v$G5_10641_out0;
assign v$RD_7489_out0 = v$G2_4640_out0;
assign v$RD_7491_out0 = v$G9_10592_out0;
assign v$RD_7493_out0 = v$G1_1929_out0;
assign v$RD_7494_out0 = v$G4_361_out0;
assign v$RD_7495_out0 = v$G6_2136_out0;
assign v$RD_7496_out0 = v$G7_11282_out0;
assign v$RD_7498_out0 = v$G8_2492_out0;
assign v$RD_7499_out0 = v$G3_261_out0;
assign v$RD_7503_out0 = v$G5_10642_out0;
assign v$RD_7504_out0 = v$G2_4641_out0;
assign v$RD_7506_out0 = v$G9_10593_out0;
assign v$RD_7508_out0 = v$G1_1930_out0;
assign v$RD_7509_out0 = v$G4_362_out0;
assign v$RD_7510_out0 = v$G6_2137_out0;
assign v$RD_7511_out0 = v$G7_11283_out0;
assign v$RD_7513_out0 = v$G8_2493_out0;
assign v$RD_7514_out0 = v$G3_262_out0;
assign v$RD_7518_out0 = v$G5_10643_out0;
assign v$RD_7519_out0 = v$G2_4642_out0;
assign v$RD_7521_out0 = v$G9_10594_out0;
assign v$RD_7523_out0 = v$G1_1931_out0;
assign v$RD_7524_out0 = v$G4_363_out0;
assign v$RD_7525_out0 = v$G6_2138_out0;
assign v$RD_7526_out0 = v$G7_11284_out0;
assign v$RD_7528_out0 = v$G8_2494_out0;
assign v$RD_7529_out0 = v$G3_263_out0;
assign v$RD_7533_out0 = v$G5_10644_out0;
assign v$RD_7534_out0 = v$G2_4643_out0;
assign v$RD_7536_out0 = v$G9_10595_out0;
assign v$RD_7538_out0 = v$G1_1932_out0;
assign v$RD_7539_out0 = v$G4_364_out0;
assign v$RD_7540_out0 = v$G6_2139_out0;
assign v$RD_7541_out0 = v$G7_11285_out0;
assign v$RD_7543_out0 = v$G8_2495_out0;
assign v$RD_7544_out0 = v$G3_264_out0;
assign v$RD_7548_out0 = v$G5_10645_out0;
assign v$RD_7549_out0 = v$G2_4644_out0;
assign v$RD_7551_out0 = v$G9_10596_out0;
assign v$RD_7553_out0 = v$G1_1933_out0;
assign v$RD_7554_out0 = v$G4_365_out0;
assign v$RD_7555_out0 = v$G6_2140_out0;
assign v$RD_7556_out0 = v$G7_11286_out0;
assign v$RD_7558_out0 = v$G8_2496_out0;
assign v$RD_7559_out0 = v$G3_265_out0;
assign v$RD_7563_out0 = v$G5_10646_out0;
assign v$RD_7564_out0 = v$G2_4645_out0;
assign v$RD_7566_out0 = v$G9_10597_out0;
assign v$RD_7568_out0 = v$G1_1934_out0;
assign v$RD_7569_out0 = v$G4_366_out0;
assign v$RD_7570_out0 = v$G6_2141_out0;
assign v$RD_7571_out0 = v$G7_11287_out0;
assign v$RD_7573_out0 = v$G8_2497_out0;
assign v$RD_7574_out0 = v$G3_266_out0;
assign v$RD_7578_out0 = v$G5_10647_out0;
assign v$RD_7579_out0 = v$G2_4646_out0;
assign v$RD_7581_out0 = v$G9_10598_out0;
assign v$RD_7583_out0 = v$G1_1935_out0;
assign v$RD_7584_out0 = v$G4_367_out0;
assign v$RD_7585_out0 = v$G6_2142_out0;
assign v$RD_7586_out0 = v$G7_11288_out0;
assign v$RD_7588_out0 = v$G8_2498_out0;
assign v$RD_7589_out0 = v$G3_267_out0;
assign v$RD_7593_out0 = v$G5_10648_out0;
assign v$RD_7594_out0 = v$G2_4647_out0;
assign v$RD_7596_out0 = v$G9_10599_out0;
assign v$RD_7598_out0 = v$G1_1936_out0;
assign v$RD_7599_out0 = v$G4_368_out0;
assign v$RD_7600_out0 = v$G6_2143_out0;
assign v$RD_7601_out0 = v$G7_11289_out0;
assign v$RD_7603_out0 = v$G8_2499_out0;
assign v$RD_7604_out0 = v$G3_268_out0;
assign v$RD_7608_out0 = v$G5_10649_out0;
assign v$RD_7609_out0 = v$G2_4648_out0;
assign v$RD_7611_out0 = v$G9_10600_out0;
assign v$RD_7613_out0 = v$G1_1937_out0;
assign v$RD_7614_out0 = v$G4_369_out0;
assign v$RD_7615_out0 = v$G6_2144_out0;
assign v$RD_7616_out0 = v$G7_11290_out0;
assign v$RD_7618_out0 = v$G8_2500_out0;
assign v$RD_7619_out0 = v$G3_269_out0;
assign v$RD_7623_out0 = v$G5_10650_out0;
assign v$RD_7624_out0 = v$G2_4649_out0;
assign v$RD_7626_out0 = v$G9_10601_out0;
assign v$RD_7628_out0 = v$G1_1938_out0;
assign v$RD_7629_out0 = v$G4_370_out0;
assign v$RD_7630_out0 = v$G6_2145_out0;
assign v$RD_7631_out0 = v$G7_11291_out0;
assign v$RD_7633_out0 = v$G8_2501_out0;
assign v$RD_7634_out0 = v$G3_270_out0;
assign v$IN_8838_out0 = v$IN_10403_out0;
assign v$IN_8839_out0 = v$IN_10404_out0;
assign v$_10372_out0 = { v$_3215_out0,v$_3278_out0 };
assign v$_10374_out0 = { v$_3217_out0,v$_3280_out0 };
assign v$_11049_out0 = v$IN_10403_out0[13:0];
assign v$_11049_out1 = v$IN_10403_out0[15:2];
assign v$_11050_out0 = v$IN_10404_out0[13:0];
assign v$_11050_out1 = v$IN_10404_out0[15:2];
assign v$G12_13221_out0 = v$RD_13567_out0 && v$_2273_out0;
assign v$G12_13224_out0 = v$RD_13570_out0 && v$_2276_out0;
assign v$G12_13226_out0 = v$RD_13572_out0 && v$_2278_out0;
assign v$G12_13227_out0 = v$RD_13573_out0 && v$_2279_out0;
assign v$G12_13228_out0 = v$RD_13574_out0 && v$_2280_out0;
assign v$G12_13229_out0 = v$RD_13575_out0 && v$_2281_out0;
assign v$G12_13230_out0 = v$RD_13576_out0 && v$_2282_out0;
assign v$G12_13231_out0 = v$RD_13577_out0 && v$_2283_out0;
assign v$G12_13232_out0 = v$RD_13578_out0 && v$_2284_out0;
assign v$G12_13233_out0 = v$RD_13579_out0 && v$_2285_out0;
assign v$G12_13234_out0 = v$RD_13580_out0 && v$_2286_out0;
assign v$G12_13235_out0 = v$RD_13581_out0 && v$_2287_out0;
assign v$G12_13236_out0 = v$RD_13582_out0 && v$_2288_out0;
assign v$G12_13239_out0 = v$RD_13585_out0 && v$_2291_out0;
assign v$G12_13241_out0 = v$RD_13587_out0 && v$_2293_out0;
assign v$G12_13242_out0 = v$RD_13588_out0 && v$_2294_out0;
assign v$G12_13243_out0 = v$RD_13589_out0 && v$_2295_out0;
assign v$G12_13244_out0 = v$RD_13590_out0 && v$_2296_out0;
assign v$G12_13245_out0 = v$RD_13591_out0 && v$_2297_out0;
assign v$G12_13246_out0 = v$RD_13592_out0 && v$_2298_out0;
assign v$G12_13247_out0 = v$RD_13593_out0 && v$_2299_out0;
assign v$G12_13248_out0 = v$RD_13594_out0 && v$_2300_out0;
assign v$G12_13249_out0 = v$RD_13595_out0 && v$_2301_out0;
assign v$G12_13250_out0 = v$RD_13596_out0 && v$_2302_out0;
assign v$G13_13352_out0 = v$RD_13567_out0 && v$_13715_out0;
assign v$G13_13355_out0 = v$RD_13570_out0 && v$_13718_out0;
assign v$G13_13357_out0 = v$RD_13572_out0 && v$_13720_out0;
assign v$G13_13358_out0 = v$RD_13573_out0 && v$_13721_out0;
assign v$G13_13359_out0 = v$RD_13574_out0 && v$_13722_out0;
assign v$G13_13360_out0 = v$RD_13575_out0 && v$_13723_out0;
assign v$G13_13361_out0 = v$RD_13576_out0 && v$_13724_out0;
assign v$G13_13362_out0 = v$RD_13577_out0 && v$_13725_out0;
assign v$G13_13363_out0 = v$RD_13578_out0 && v$_13726_out0;
assign v$G13_13364_out0 = v$RD_13579_out0 && v$_13727_out0;
assign v$G13_13365_out0 = v$RD_13580_out0 && v$_13728_out0;
assign v$G13_13366_out0 = v$RD_13581_out0 && v$_13729_out0;
assign v$G13_13367_out0 = v$RD_13582_out0 && v$_13730_out0;
assign v$G13_13370_out0 = v$RD_13585_out0 && v$_13733_out0;
assign v$G13_13372_out0 = v$RD_13587_out0 && v$_13735_out0;
assign v$G13_13373_out0 = v$RD_13588_out0 && v$_13736_out0;
assign v$G13_13374_out0 = v$RD_13589_out0 && v$_13737_out0;
assign v$G13_13375_out0 = v$RD_13590_out0 && v$_13738_out0;
assign v$G13_13376_out0 = v$RD_13591_out0 && v$_13739_out0;
assign v$G13_13377_out0 = v$RD_13592_out0 && v$_13740_out0;
assign v$G13_13378_out0 = v$RD_13593_out0 && v$_13741_out0;
assign v$G13_13379_out0 = v$RD_13594_out0 && v$_13742_out0;
assign v$G13_13380_out0 = v$RD_13595_out0 && v$_13743_out0;
assign v$G13_13381_out0 = v$RD_13596_out0 && v$_13744_out0;
assign v$IN_13668_out0 = v$SIG$TO$SHIFT_5836_out0;
assign v$IN_13669_out0 = v$SIG$TO$SHIFT_5837_out0;
assign v$G14_13672_out0 = v$RD_13567_out0 && v$_6830_out0;
assign v$G14_13675_out0 = v$RD_13570_out0 && v$_6833_out0;
assign v$G14_13677_out0 = v$RD_13572_out0 && v$_6835_out0;
assign v$G14_13678_out0 = v$RD_13573_out0 && v$_6836_out0;
assign v$G14_13679_out0 = v$RD_13574_out0 && v$_6837_out0;
assign v$G14_13680_out0 = v$RD_13575_out0 && v$_6838_out0;
assign v$G14_13681_out0 = v$RD_13576_out0 && v$_6839_out0;
assign v$G14_13682_out0 = v$RD_13577_out0 && v$_6840_out0;
assign v$G14_13683_out0 = v$RD_13578_out0 && v$_6841_out0;
assign v$G14_13684_out0 = v$RD_13579_out0 && v$_6842_out0;
assign v$G14_13685_out0 = v$RD_13580_out0 && v$_6843_out0;
assign v$G14_13686_out0 = v$RD_13581_out0 && v$_6844_out0;
assign v$G14_13687_out0 = v$RD_13582_out0 && v$_6845_out0;
assign v$G14_13690_out0 = v$RD_13585_out0 && v$_6848_out0;
assign v$G14_13692_out0 = v$RD_13587_out0 && v$_6850_out0;
assign v$G14_13693_out0 = v$RD_13588_out0 && v$_6851_out0;
assign v$G14_13694_out0 = v$RD_13589_out0 && v$_6852_out0;
assign v$G14_13695_out0 = v$RD_13590_out0 && v$_6853_out0;
assign v$G14_13696_out0 = v$RD_13591_out0 && v$_6854_out0;
assign v$G14_13697_out0 = v$RD_13592_out0 && v$_6855_out0;
assign v$G14_13698_out0 = v$RD_13593_out0 && v$_6856_out0;
assign v$G14_13699_out0 = v$RD_13594_out0 && v$_6857_out0;
assign v$G14_13700_out0 = v$RD_13595_out0 && v$_6858_out0;
assign v$G14_13701_out0 = v$RD_13596_out0 && v$_6859_out0;
assign v$IN1_2189_out0 = v$IN_13668_out0;
assign v$IN1_2190_out0 = v$IN_13669_out0;
assign v$NOTUSED_2589_out0 = v$_11049_out1;
assign v$NOTUSED_2590_out0 = v$_11050_out1;
assign v$_2684_out0 = { v$_10372_out0,v$_113_out0 };
assign v$_2686_out0 = { v$_10374_out0,v$_115_out0 };
assign v$_4449_out0 = { v$_2345_out0,v$_449_out0 };
assign v$_4451_out0 = { v$_2347_out0,v$_451_out0 };
assign v$RD_5868_out0 = v$RD_7190_out0;
assign v$RD_5870_out0 = v$RD_7191_out0;
assign v$RD_5875_out0 = v$RD_7193_out0;
assign v$RD_5879_out0 = v$RD_7195_out0;
assign v$RD_5881_out0 = v$RD_7196_out0;
assign v$RD_5883_out0 = v$RD_7197_out0;
assign v$RD_5885_out0 = v$RD_7198_out0;
assign v$RD_5889_out0 = v$RD_7200_out0;
assign v$RD_5891_out0 = v$RD_7201_out0;
assign v$RD_5893_out0 = v$RD_7202_out0;
assign v$RD_5895_out0 = v$RD_7203_out0;
assign v$RD_5901_out0 = v$RD_7206_out0;
assign v$RD_5907_out0 = v$RD_7208_out0;
assign v$RD_5917_out0 = v$RD_7213_out0;
assign v$RD_5923_out0 = v$RD_7216_out0;
assign v$RD_5925_out0 = v$RD_7217_out0;
assign v$RD_5927_out0 = v$RD_7218_out0;
assign v$RD_5933_out0 = v$RD_7221_out0;
assign v$RD_5938_out0 = v$RD_7223_out0;
assign v$RD_5948_out0 = v$RD_7228_out0;
assign v$RD_5960_out0 = v$RD_7234_out0;
assign v$RD_5962_out0 = v$RD_7235_out0;
assign v$RD_5967_out0 = v$RD_7237_out0;
assign v$RD_5971_out0 = v$RD_7239_out0;
assign v$RD_5973_out0 = v$RD_7240_out0;
assign v$RD_5975_out0 = v$RD_7241_out0;
assign v$RD_5977_out0 = v$RD_7242_out0;
assign v$RD_5981_out0 = v$RD_7244_out0;
assign v$RD_5983_out0 = v$RD_7245_out0;
assign v$RD_5985_out0 = v$RD_7246_out0;
assign v$RD_5987_out0 = v$RD_7247_out0;
assign v$RD_5989_out0 = v$RD_7248_out0;
assign v$RD_5995_out0 = v$RD_7251_out0;
assign v$RD_6000_out0 = v$RD_7253_out0;
assign v$RD_6010_out0 = v$RD_7258_out0;
assign v$RD_6022_out0 = v$RD_7264_out0;
assign v$RD_6024_out0 = v$RD_7265_out0;
assign v$RD_6029_out0 = v$RD_7267_out0;
assign v$RD_6033_out0 = v$RD_7269_out0;
assign v$RD_6035_out0 = v$RD_7270_out0;
assign v$RD_6037_out0 = v$RD_7271_out0;
assign v$RD_6039_out0 = v$RD_7272_out0;
assign v$RD_6043_out0 = v$RD_7274_out0;
assign v$RD_6045_out0 = v$RD_7275_out0;
assign v$RD_6053_out0 = v$RD_7279_out0;
assign v$RD_6055_out0 = v$RD_7280_out0;
assign v$RD_6060_out0 = v$RD_7282_out0;
assign v$RD_6064_out0 = v$RD_7284_out0;
assign v$RD_6066_out0 = v$RD_7285_out0;
assign v$RD_6068_out0 = v$RD_7286_out0;
assign v$RD_6070_out0 = v$RD_7287_out0;
assign v$RD_6074_out0 = v$RD_7289_out0;
assign v$RD_6076_out0 = v$RD_7290_out0;
assign v$RD_6084_out0 = v$RD_7294_out0;
assign v$RD_6086_out0 = v$RD_7295_out0;
assign v$RD_6091_out0 = v$RD_7297_out0;
assign v$RD_6095_out0 = v$RD_7299_out0;
assign v$RD_6097_out0 = v$RD_7300_out0;
assign v$RD_6099_out0 = v$RD_7301_out0;
assign v$RD_6101_out0 = v$RD_7302_out0;
assign v$RD_6105_out0 = v$RD_7304_out0;
assign v$RD_6107_out0 = v$RD_7305_out0;
assign v$RD_6115_out0 = v$RD_7309_out0;
assign v$RD_6117_out0 = v$RD_7310_out0;
assign v$RD_6122_out0 = v$RD_7312_out0;
assign v$RD_6126_out0 = v$RD_7314_out0;
assign v$RD_6128_out0 = v$RD_7315_out0;
assign v$RD_6130_out0 = v$RD_7316_out0;
assign v$RD_6132_out0 = v$RD_7317_out0;
assign v$RD_6136_out0 = v$RD_7319_out0;
assign v$RD_6138_out0 = v$RD_7320_out0;
assign v$RD_6146_out0 = v$RD_7324_out0;
assign v$RD_6148_out0 = v$RD_7325_out0;
assign v$RD_6153_out0 = v$RD_7327_out0;
assign v$RD_6157_out0 = v$RD_7329_out0;
assign v$RD_6159_out0 = v$RD_7330_out0;
assign v$RD_6161_out0 = v$RD_7331_out0;
assign v$RD_6163_out0 = v$RD_7332_out0;
assign v$RD_6167_out0 = v$RD_7334_out0;
assign v$RD_6169_out0 = v$RD_7335_out0;
assign v$RD_6177_out0 = v$RD_7339_out0;
assign v$RD_6179_out0 = v$RD_7340_out0;
assign v$RD_6184_out0 = v$RD_7342_out0;
assign v$RD_6188_out0 = v$RD_7344_out0;
assign v$RD_6190_out0 = v$RD_7345_out0;
assign v$RD_6192_out0 = v$RD_7346_out0;
assign v$RD_6194_out0 = v$RD_7347_out0;
assign v$RD_6198_out0 = v$RD_7349_out0;
assign v$RD_6200_out0 = v$RD_7350_out0;
assign v$RD_6208_out0 = v$RD_7354_out0;
assign v$RD_6210_out0 = v$RD_7355_out0;
assign v$RD_6215_out0 = v$RD_7357_out0;
assign v$RD_6219_out0 = v$RD_7359_out0;
assign v$RD_6221_out0 = v$RD_7360_out0;
assign v$RD_6223_out0 = v$RD_7361_out0;
assign v$RD_6225_out0 = v$RD_7362_out0;
assign v$RD_6229_out0 = v$RD_7364_out0;
assign v$RD_6231_out0 = v$RD_7365_out0;
assign v$RD_6239_out0 = v$RD_7369_out0;
assign v$RD_6241_out0 = v$RD_7370_out0;
assign v$RD_6246_out0 = v$RD_7372_out0;
assign v$RD_6250_out0 = v$RD_7374_out0;
assign v$RD_6252_out0 = v$RD_7375_out0;
assign v$RD_6254_out0 = v$RD_7376_out0;
assign v$RD_6256_out0 = v$RD_7377_out0;
assign v$RD_6260_out0 = v$RD_7379_out0;
assign v$RD_6262_out0 = v$RD_7380_out0;
assign v$RD_6270_out0 = v$RD_7384_out0;
assign v$RD_6272_out0 = v$RD_7385_out0;
assign v$RD_6277_out0 = v$RD_7387_out0;
assign v$RD_6281_out0 = v$RD_7389_out0;
assign v$RD_6283_out0 = v$RD_7390_out0;
assign v$RD_6285_out0 = v$RD_7391_out0;
assign v$RD_6287_out0 = v$RD_7392_out0;
assign v$RD_6291_out0 = v$RD_7394_out0;
assign v$RD_6293_out0 = v$RD_7395_out0;
assign v$RD_6301_out0 = v$RD_7399_out0;
assign v$RD_6303_out0 = v$RD_7400_out0;
assign v$RD_6308_out0 = v$RD_7402_out0;
assign v$RD_6312_out0 = v$RD_7404_out0;
assign v$RD_6314_out0 = v$RD_7405_out0;
assign v$RD_6316_out0 = v$RD_7406_out0;
assign v$RD_6318_out0 = v$RD_7407_out0;
assign v$RD_6322_out0 = v$RD_7409_out0;
assign v$RD_6324_out0 = v$RD_7410_out0;
assign v$RD_6332_out0 = v$RD_7414_out0;
assign v$RD_6334_out0 = v$RD_7415_out0;
assign v$RD_6339_out0 = v$RD_7417_out0;
assign v$RD_6343_out0 = v$RD_7419_out0;
assign v$RD_6345_out0 = v$RD_7420_out0;
assign v$RD_6347_out0 = v$RD_7421_out0;
assign v$RD_6349_out0 = v$RD_7422_out0;
assign v$RD_6353_out0 = v$RD_7424_out0;
assign v$RD_6355_out0 = v$RD_7425_out0;
assign v$RD_6357_out0 = v$RD_7426_out0;
assign v$RD_6359_out0 = v$RD_7427_out0;
assign v$RD_6365_out0 = v$RD_7430_out0;
assign v$RD_6371_out0 = v$RD_7432_out0;
assign v$RD_6381_out0 = v$RD_7437_out0;
assign v$RD_6387_out0 = v$RD_7440_out0;
assign v$RD_6389_out0 = v$RD_7441_out0;
assign v$RD_6391_out0 = v$RD_7442_out0;
assign v$RD_6397_out0 = v$RD_7445_out0;
assign v$RD_6402_out0 = v$RD_7447_out0;
assign v$RD_6412_out0 = v$RD_7452_out0;
assign v$RD_6424_out0 = v$RD_7458_out0;
assign v$RD_6426_out0 = v$RD_7459_out0;
assign v$RD_6431_out0 = v$RD_7461_out0;
assign v$RD_6435_out0 = v$RD_7463_out0;
assign v$RD_6437_out0 = v$RD_7464_out0;
assign v$RD_6439_out0 = v$RD_7465_out0;
assign v$RD_6441_out0 = v$RD_7466_out0;
assign v$RD_6445_out0 = v$RD_7468_out0;
assign v$RD_6447_out0 = v$RD_7469_out0;
assign v$RD_6449_out0 = v$RD_7470_out0;
assign v$RD_6451_out0 = v$RD_7471_out0;
assign v$RD_6453_out0 = v$RD_7472_out0;
assign v$RD_6459_out0 = v$RD_7475_out0;
assign v$RD_6464_out0 = v$RD_7477_out0;
assign v$RD_6474_out0 = v$RD_7482_out0;
assign v$RD_6486_out0 = v$RD_7488_out0;
assign v$RD_6488_out0 = v$RD_7489_out0;
assign v$RD_6493_out0 = v$RD_7491_out0;
assign v$RD_6497_out0 = v$RD_7493_out0;
assign v$RD_6499_out0 = v$RD_7494_out0;
assign v$RD_6501_out0 = v$RD_7495_out0;
assign v$RD_6503_out0 = v$RD_7496_out0;
assign v$RD_6507_out0 = v$RD_7498_out0;
assign v$RD_6509_out0 = v$RD_7499_out0;
assign v$RD_6517_out0 = v$RD_7503_out0;
assign v$RD_6519_out0 = v$RD_7504_out0;
assign v$RD_6524_out0 = v$RD_7506_out0;
assign v$RD_6528_out0 = v$RD_7508_out0;
assign v$RD_6530_out0 = v$RD_7509_out0;
assign v$RD_6532_out0 = v$RD_7510_out0;
assign v$RD_6534_out0 = v$RD_7511_out0;
assign v$RD_6538_out0 = v$RD_7513_out0;
assign v$RD_6540_out0 = v$RD_7514_out0;
assign v$RD_6548_out0 = v$RD_7518_out0;
assign v$RD_6550_out0 = v$RD_7519_out0;
assign v$RD_6555_out0 = v$RD_7521_out0;
assign v$RD_6559_out0 = v$RD_7523_out0;
assign v$RD_6561_out0 = v$RD_7524_out0;
assign v$RD_6563_out0 = v$RD_7525_out0;
assign v$RD_6565_out0 = v$RD_7526_out0;
assign v$RD_6569_out0 = v$RD_7528_out0;
assign v$RD_6571_out0 = v$RD_7529_out0;
assign v$RD_6579_out0 = v$RD_7533_out0;
assign v$RD_6581_out0 = v$RD_7534_out0;
assign v$RD_6586_out0 = v$RD_7536_out0;
assign v$RD_6590_out0 = v$RD_7538_out0;
assign v$RD_6592_out0 = v$RD_7539_out0;
assign v$RD_6594_out0 = v$RD_7540_out0;
assign v$RD_6596_out0 = v$RD_7541_out0;
assign v$RD_6600_out0 = v$RD_7543_out0;
assign v$RD_6602_out0 = v$RD_7544_out0;
assign v$RD_6610_out0 = v$RD_7548_out0;
assign v$RD_6612_out0 = v$RD_7549_out0;
assign v$RD_6617_out0 = v$RD_7551_out0;
assign v$RD_6621_out0 = v$RD_7553_out0;
assign v$RD_6623_out0 = v$RD_7554_out0;
assign v$RD_6625_out0 = v$RD_7555_out0;
assign v$RD_6627_out0 = v$RD_7556_out0;
assign v$RD_6631_out0 = v$RD_7558_out0;
assign v$RD_6633_out0 = v$RD_7559_out0;
assign v$RD_6641_out0 = v$RD_7563_out0;
assign v$RD_6643_out0 = v$RD_7564_out0;
assign v$RD_6648_out0 = v$RD_7566_out0;
assign v$RD_6652_out0 = v$RD_7568_out0;
assign v$RD_6654_out0 = v$RD_7569_out0;
assign v$RD_6656_out0 = v$RD_7570_out0;
assign v$RD_6658_out0 = v$RD_7571_out0;
assign v$RD_6662_out0 = v$RD_7573_out0;
assign v$RD_6664_out0 = v$RD_7574_out0;
assign v$RD_6672_out0 = v$RD_7578_out0;
assign v$RD_6674_out0 = v$RD_7579_out0;
assign v$RD_6679_out0 = v$RD_7581_out0;
assign v$RD_6683_out0 = v$RD_7583_out0;
assign v$RD_6685_out0 = v$RD_7584_out0;
assign v$RD_6687_out0 = v$RD_7585_out0;
assign v$RD_6689_out0 = v$RD_7586_out0;
assign v$RD_6693_out0 = v$RD_7588_out0;
assign v$RD_6695_out0 = v$RD_7589_out0;
assign v$RD_6703_out0 = v$RD_7593_out0;
assign v$RD_6705_out0 = v$RD_7594_out0;
assign v$RD_6710_out0 = v$RD_7596_out0;
assign v$RD_6714_out0 = v$RD_7598_out0;
assign v$RD_6716_out0 = v$RD_7599_out0;
assign v$RD_6718_out0 = v$RD_7600_out0;
assign v$RD_6720_out0 = v$RD_7601_out0;
assign v$RD_6724_out0 = v$RD_7603_out0;
assign v$RD_6726_out0 = v$RD_7604_out0;
assign v$RD_6734_out0 = v$RD_7608_out0;
assign v$RD_6736_out0 = v$RD_7609_out0;
assign v$RD_6741_out0 = v$RD_7611_out0;
assign v$RD_6745_out0 = v$RD_7613_out0;
assign v$RD_6747_out0 = v$RD_7614_out0;
assign v$RD_6749_out0 = v$RD_7615_out0;
assign v$RD_6751_out0 = v$RD_7616_out0;
assign v$RD_6755_out0 = v$RD_7618_out0;
assign v$RD_6757_out0 = v$RD_7619_out0;
assign v$RD_6765_out0 = v$RD_7623_out0;
assign v$RD_6767_out0 = v$RD_7624_out0;
assign v$RD_6772_out0 = v$RD_7626_out0;
assign v$RD_6776_out0 = v$RD_7628_out0;
assign v$RD_6778_out0 = v$RD_7629_out0;
assign v$RD_6780_out0 = v$RD_7630_out0;
assign v$RD_6782_out0 = v$RD_7631_out0;
assign v$RD_6786_out0 = v$RD_7633_out0;
assign v$RD_6788_out0 = v$RD_7634_out0;
assign v$RD_7187_out0 = v$G12_13221_out0;
assign v$RD_7188_out0 = v$G14_13672_out0;
assign v$RD_7189_out0 = v$G15_132_out0;
assign v$RD_7192_out0 = v$G13_13352_out0;
assign v$RD_7194_out0 = v$G10_6975_out0;
assign v$RD_7199_out0 = v$G11_651_out0;
assign v$RD_7231_out0 = v$G12_13224_out0;
assign v$RD_7232_out0 = v$G14_13675_out0;
assign v$RD_7233_out0 = v$G15_135_out0;
assign v$RD_7236_out0 = v$G13_13355_out0;
assign v$RD_7238_out0 = v$G10_6978_out0;
assign v$RD_7243_out0 = v$G11_654_out0;
assign v$RD_7261_out0 = v$G12_13226_out0;
assign v$RD_7262_out0 = v$G14_13677_out0;
assign v$RD_7263_out0 = v$G15_137_out0;
assign v$RD_7266_out0 = v$G13_13357_out0;
assign v$RD_7268_out0 = v$G10_6980_out0;
assign v$RD_7273_out0 = v$G11_656_out0;
assign v$RD_7276_out0 = v$G12_13227_out0;
assign v$RD_7277_out0 = v$G14_13678_out0;
assign v$RD_7278_out0 = v$G15_138_out0;
assign v$RD_7281_out0 = v$G13_13358_out0;
assign v$RD_7283_out0 = v$G10_6981_out0;
assign v$RD_7288_out0 = v$G11_657_out0;
assign v$RD_7291_out0 = v$G12_13228_out0;
assign v$RD_7292_out0 = v$G14_13679_out0;
assign v$RD_7293_out0 = v$G15_139_out0;
assign v$RD_7296_out0 = v$G13_13359_out0;
assign v$RD_7298_out0 = v$G10_6982_out0;
assign v$RD_7303_out0 = v$G11_658_out0;
assign v$RD_7306_out0 = v$G12_13229_out0;
assign v$RD_7307_out0 = v$G14_13680_out0;
assign v$RD_7308_out0 = v$G15_140_out0;
assign v$RD_7311_out0 = v$G13_13360_out0;
assign v$RD_7313_out0 = v$G10_6983_out0;
assign v$RD_7318_out0 = v$G11_659_out0;
assign v$RD_7321_out0 = v$G12_13230_out0;
assign v$RD_7322_out0 = v$G14_13681_out0;
assign v$RD_7323_out0 = v$G15_141_out0;
assign v$RD_7326_out0 = v$G13_13361_out0;
assign v$RD_7328_out0 = v$G10_6984_out0;
assign v$RD_7333_out0 = v$G11_660_out0;
assign v$RD_7336_out0 = v$G12_13231_out0;
assign v$RD_7337_out0 = v$G14_13682_out0;
assign v$RD_7338_out0 = v$G15_142_out0;
assign v$RD_7341_out0 = v$G13_13362_out0;
assign v$RD_7343_out0 = v$G10_6985_out0;
assign v$RD_7348_out0 = v$G11_661_out0;
assign v$RD_7351_out0 = v$G12_13232_out0;
assign v$RD_7352_out0 = v$G14_13683_out0;
assign v$RD_7353_out0 = v$G15_143_out0;
assign v$RD_7356_out0 = v$G13_13363_out0;
assign v$RD_7358_out0 = v$G10_6986_out0;
assign v$RD_7363_out0 = v$G11_662_out0;
assign v$RD_7366_out0 = v$G12_13233_out0;
assign v$RD_7367_out0 = v$G14_13684_out0;
assign v$RD_7368_out0 = v$G15_144_out0;
assign v$RD_7371_out0 = v$G13_13364_out0;
assign v$RD_7373_out0 = v$G10_6987_out0;
assign v$RD_7378_out0 = v$G11_663_out0;
assign v$RD_7381_out0 = v$G12_13234_out0;
assign v$RD_7382_out0 = v$G14_13685_out0;
assign v$RD_7383_out0 = v$G15_145_out0;
assign v$RD_7386_out0 = v$G13_13365_out0;
assign v$RD_7388_out0 = v$G10_6988_out0;
assign v$RD_7393_out0 = v$G11_664_out0;
assign v$RD_7396_out0 = v$G12_13235_out0;
assign v$RD_7397_out0 = v$G14_13686_out0;
assign v$RD_7398_out0 = v$G15_146_out0;
assign v$RD_7401_out0 = v$G13_13366_out0;
assign v$RD_7403_out0 = v$G10_6989_out0;
assign v$RD_7408_out0 = v$G11_665_out0;
assign v$RD_7411_out0 = v$G12_13236_out0;
assign v$RD_7412_out0 = v$G14_13687_out0;
assign v$RD_7413_out0 = v$G15_147_out0;
assign v$RD_7416_out0 = v$G13_13367_out0;
assign v$RD_7418_out0 = v$G10_6990_out0;
assign v$RD_7423_out0 = v$G11_666_out0;
assign v$RD_7455_out0 = v$G12_13239_out0;
assign v$RD_7456_out0 = v$G14_13690_out0;
assign v$RD_7457_out0 = v$G15_150_out0;
assign v$RD_7460_out0 = v$G13_13370_out0;
assign v$RD_7462_out0 = v$G10_6993_out0;
assign v$RD_7467_out0 = v$G11_669_out0;
assign v$RD_7485_out0 = v$G12_13241_out0;
assign v$RD_7486_out0 = v$G14_13692_out0;
assign v$RD_7487_out0 = v$G15_152_out0;
assign v$RD_7490_out0 = v$G13_13372_out0;
assign v$RD_7492_out0 = v$G10_6995_out0;
assign v$RD_7497_out0 = v$G11_671_out0;
assign v$RD_7500_out0 = v$G12_13242_out0;
assign v$RD_7501_out0 = v$G14_13693_out0;
assign v$RD_7502_out0 = v$G15_153_out0;
assign v$RD_7505_out0 = v$G13_13373_out0;
assign v$RD_7507_out0 = v$G10_6996_out0;
assign v$RD_7512_out0 = v$G11_672_out0;
assign v$RD_7515_out0 = v$G12_13243_out0;
assign v$RD_7516_out0 = v$G14_13694_out0;
assign v$RD_7517_out0 = v$G15_154_out0;
assign v$RD_7520_out0 = v$G13_13374_out0;
assign v$RD_7522_out0 = v$G10_6997_out0;
assign v$RD_7527_out0 = v$G11_673_out0;
assign v$RD_7530_out0 = v$G12_13244_out0;
assign v$RD_7531_out0 = v$G14_13695_out0;
assign v$RD_7532_out0 = v$G15_155_out0;
assign v$RD_7535_out0 = v$G13_13375_out0;
assign v$RD_7537_out0 = v$G10_6998_out0;
assign v$RD_7542_out0 = v$G11_674_out0;
assign v$RD_7545_out0 = v$G12_13245_out0;
assign v$RD_7546_out0 = v$G14_13696_out0;
assign v$RD_7547_out0 = v$G15_156_out0;
assign v$RD_7550_out0 = v$G13_13376_out0;
assign v$RD_7552_out0 = v$G10_6999_out0;
assign v$RD_7557_out0 = v$G11_675_out0;
assign v$RD_7560_out0 = v$G12_13246_out0;
assign v$RD_7561_out0 = v$G14_13697_out0;
assign v$RD_7562_out0 = v$G15_157_out0;
assign v$RD_7565_out0 = v$G13_13377_out0;
assign v$RD_7567_out0 = v$G10_7000_out0;
assign v$RD_7572_out0 = v$G11_676_out0;
assign v$RD_7575_out0 = v$G12_13247_out0;
assign v$RD_7576_out0 = v$G14_13698_out0;
assign v$RD_7577_out0 = v$G15_158_out0;
assign v$RD_7580_out0 = v$G13_13378_out0;
assign v$RD_7582_out0 = v$G10_7001_out0;
assign v$RD_7587_out0 = v$G11_677_out0;
assign v$RD_7590_out0 = v$G12_13248_out0;
assign v$RD_7591_out0 = v$G14_13699_out0;
assign v$RD_7592_out0 = v$G15_159_out0;
assign v$RD_7595_out0 = v$G13_13379_out0;
assign v$RD_7597_out0 = v$G10_7002_out0;
assign v$RD_7602_out0 = v$G11_678_out0;
assign v$RD_7605_out0 = v$G12_13249_out0;
assign v$RD_7606_out0 = v$G14_13700_out0;
assign v$RD_7607_out0 = v$G15_160_out0;
assign v$RD_7610_out0 = v$G13_13380_out0;
assign v$RD_7612_out0 = v$G10_7003_out0;
assign v$RD_7617_out0 = v$G11_679_out0;
assign v$RD_7620_out0 = v$G12_13250_out0;
assign v$RD_7621_out0 = v$G14_13701_out0;
assign v$RD_7622_out0 = v$G15_161_out0;
assign v$RD_7625_out0 = v$G13_13381_out0;
assign v$RD_7627_out0 = v$G10_7004_out0;
assign v$RD_7632_out0 = v$G11_680_out0;
assign v$ADDER$IN_8745_out0 = v$_1212_out0;
assign v$ADDER$IN_8747_out0 = v$_1214_out0;
assign v$_10333_out0 = { v$C1_11292_out0,v$_11049_out0 };
assign v$_10334_out0 = { v$C1_11293_out0,v$_11050_out0 };
assign v$_10783_out0 = { v$_4733_out0,v$G12_4699_out0 };
assign v$MUX1_6_out0 = v$LSL_2842_out0 ? v$_10333_out0 : v$IN_8838_out0;
assign v$MUX1_7_out0 = v$LSL_2843_out0 ? v$_10334_out0 : v$IN_8839_out0;
assign v$_1867_out0 = { v$_2684_out0,v$_4449_out0 };
assign v$_1869_out0 = { v$_2686_out0,v$_4451_out0 };
assign {v$A1_3174_out1,v$A1_3174_out0 } = v$RM_13508_out0 + v$ADDER$IN_8745_out0 + v$U_10469_out0;
assign {v$A1_3175_out1,v$A1_3175_out0 } = v$RM_13509_out0 + v$ADDER$IN_8747_out0 + v$U_10470_out0;
assign v$_3907_out0 = v$IN1_2189_out0[0:0];
assign v$_3907_out1 = v$IN1_2189_out0[10:10];
assign v$_3908_out0 = v$IN1_2190_out0[0:0];
assign v$_3908_out1 = v$IN1_2190_out0[10:10];
assign v$RD_5862_out0 = v$RD_7187_out0;
assign v$RD_5864_out0 = v$RD_7188_out0;
assign v$RD_5866_out0 = v$RD_7189_out0;
assign v$RD_5872_out0 = v$RD_7192_out0;
assign v$RD_5877_out0 = v$RD_7194_out0;
assign v$RD_5887_out0 = v$RD_7199_out0;
assign v$RD_5954_out0 = v$RD_7231_out0;
assign v$RD_5956_out0 = v$RD_7232_out0;
assign v$RD_5958_out0 = v$RD_7233_out0;
assign v$RD_5964_out0 = v$RD_7236_out0;
assign v$RD_5969_out0 = v$RD_7238_out0;
assign v$RD_5979_out0 = v$RD_7243_out0;
assign v$RD_6016_out0 = v$RD_7261_out0;
assign v$RD_6018_out0 = v$RD_7262_out0;
assign v$RD_6020_out0 = v$RD_7263_out0;
assign v$RD_6026_out0 = v$RD_7266_out0;
assign v$RD_6031_out0 = v$RD_7268_out0;
assign v$RD_6041_out0 = v$RD_7273_out0;
assign v$RD_6047_out0 = v$RD_7276_out0;
assign v$RD_6049_out0 = v$RD_7277_out0;
assign v$RD_6051_out0 = v$RD_7278_out0;
assign v$RD_6057_out0 = v$RD_7281_out0;
assign v$RD_6062_out0 = v$RD_7283_out0;
assign v$RD_6072_out0 = v$RD_7288_out0;
assign v$RD_6078_out0 = v$RD_7291_out0;
assign v$RD_6080_out0 = v$RD_7292_out0;
assign v$RD_6082_out0 = v$RD_7293_out0;
assign v$RD_6088_out0 = v$RD_7296_out0;
assign v$RD_6093_out0 = v$RD_7298_out0;
assign v$RD_6103_out0 = v$RD_7303_out0;
assign v$RD_6109_out0 = v$RD_7306_out0;
assign v$RD_6111_out0 = v$RD_7307_out0;
assign v$RD_6113_out0 = v$RD_7308_out0;
assign v$RD_6119_out0 = v$RD_7311_out0;
assign v$RD_6124_out0 = v$RD_7313_out0;
assign v$RD_6134_out0 = v$RD_7318_out0;
assign v$RD_6140_out0 = v$RD_7321_out0;
assign v$RD_6142_out0 = v$RD_7322_out0;
assign v$RD_6144_out0 = v$RD_7323_out0;
assign v$RD_6150_out0 = v$RD_7326_out0;
assign v$RD_6155_out0 = v$RD_7328_out0;
assign v$RD_6165_out0 = v$RD_7333_out0;
assign v$RD_6171_out0 = v$RD_7336_out0;
assign v$RD_6173_out0 = v$RD_7337_out0;
assign v$RD_6175_out0 = v$RD_7338_out0;
assign v$RD_6181_out0 = v$RD_7341_out0;
assign v$RD_6186_out0 = v$RD_7343_out0;
assign v$RD_6196_out0 = v$RD_7348_out0;
assign v$RD_6202_out0 = v$RD_7351_out0;
assign v$RD_6204_out0 = v$RD_7352_out0;
assign v$RD_6206_out0 = v$RD_7353_out0;
assign v$RD_6212_out0 = v$RD_7356_out0;
assign v$RD_6217_out0 = v$RD_7358_out0;
assign v$RD_6227_out0 = v$RD_7363_out0;
assign v$RD_6233_out0 = v$RD_7366_out0;
assign v$RD_6235_out0 = v$RD_7367_out0;
assign v$RD_6237_out0 = v$RD_7368_out0;
assign v$RD_6243_out0 = v$RD_7371_out0;
assign v$RD_6248_out0 = v$RD_7373_out0;
assign v$RD_6258_out0 = v$RD_7378_out0;
assign v$RD_6264_out0 = v$RD_7381_out0;
assign v$RD_6266_out0 = v$RD_7382_out0;
assign v$RD_6268_out0 = v$RD_7383_out0;
assign v$RD_6274_out0 = v$RD_7386_out0;
assign v$RD_6279_out0 = v$RD_7388_out0;
assign v$RD_6289_out0 = v$RD_7393_out0;
assign v$RD_6295_out0 = v$RD_7396_out0;
assign v$RD_6297_out0 = v$RD_7397_out0;
assign v$RD_6299_out0 = v$RD_7398_out0;
assign v$RD_6305_out0 = v$RD_7401_out0;
assign v$RD_6310_out0 = v$RD_7403_out0;
assign v$RD_6320_out0 = v$RD_7408_out0;
assign v$RD_6326_out0 = v$RD_7411_out0;
assign v$RD_6328_out0 = v$RD_7412_out0;
assign v$RD_6330_out0 = v$RD_7413_out0;
assign v$RD_6336_out0 = v$RD_7416_out0;
assign v$RD_6341_out0 = v$RD_7418_out0;
assign v$RD_6351_out0 = v$RD_7423_out0;
assign v$RD_6418_out0 = v$RD_7455_out0;
assign v$RD_6420_out0 = v$RD_7456_out0;
assign v$RD_6422_out0 = v$RD_7457_out0;
assign v$RD_6428_out0 = v$RD_7460_out0;
assign v$RD_6433_out0 = v$RD_7462_out0;
assign v$RD_6443_out0 = v$RD_7467_out0;
assign v$RD_6480_out0 = v$RD_7485_out0;
assign v$RD_6482_out0 = v$RD_7486_out0;
assign v$RD_6484_out0 = v$RD_7487_out0;
assign v$RD_6490_out0 = v$RD_7490_out0;
assign v$RD_6495_out0 = v$RD_7492_out0;
assign v$RD_6505_out0 = v$RD_7497_out0;
assign v$RD_6511_out0 = v$RD_7500_out0;
assign v$RD_6513_out0 = v$RD_7501_out0;
assign v$RD_6515_out0 = v$RD_7502_out0;
assign v$RD_6521_out0 = v$RD_7505_out0;
assign v$RD_6526_out0 = v$RD_7507_out0;
assign v$RD_6536_out0 = v$RD_7512_out0;
assign v$RD_6542_out0 = v$RD_7515_out0;
assign v$RD_6544_out0 = v$RD_7516_out0;
assign v$RD_6546_out0 = v$RD_7517_out0;
assign v$RD_6552_out0 = v$RD_7520_out0;
assign v$RD_6557_out0 = v$RD_7522_out0;
assign v$RD_6567_out0 = v$RD_7527_out0;
assign v$RD_6573_out0 = v$RD_7530_out0;
assign v$RD_6575_out0 = v$RD_7531_out0;
assign v$RD_6577_out0 = v$RD_7532_out0;
assign v$RD_6583_out0 = v$RD_7535_out0;
assign v$RD_6588_out0 = v$RD_7537_out0;
assign v$RD_6598_out0 = v$RD_7542_out0;
assign v$RD_6604_out0 = v$RD_7545_out0;
assign v$RD_6606_out0 = v$RD_7546_out0;
assign v$RD_6608_out0 = v$RD_7547_out0;
assign v$RD_6614_out0 = v$RD_7550_out0;
assign v$RD_6619_out0 = v$RD_7552_out0;
assign v$RD_6629_out0 = v$RD_7557_out0;
assign v$RD_6635_out0 = v$RD_7560_out0;
assign v$RD_6637_out0 = v$RD_7561_out0;
assign v$RD_6639_out0 = v$RD_7562_out0;
assign v$RD_6645_out0 = v$RD_7565_out0;
assign v$RD_6650_out0 = v$RD_7567_out0;
assign v$RD_6660_out0 = v$RD_7572_out0;
assign v$RD_6666_out0 = v$RD_7575_out0;
assign v$RD_6668_out0 = v$RD_7576_out0;
assign v$RD_6670_out0 = v$RD_7577_out0;
assign v$RD_6676_out0 = v$RD_7580_out0;
assign v$RD_6681_out0 = v$RD_7582_out0;
assign v$RD_6691_out0 = v$RD_7587_out0;
assign v$RD_6697_out0 = v$RD_7590_out0;
assign v$RD_6699_out0 = v$RD_7591_out0;
assign v$RD_6701_out0 = v$RD_7592_out0;
assign v$RD_6707_out0 = v$RD_7595_out0;
assign v$RD_6712_out0 = v$RD_7597_out0;
assign v$RD_6722_out0 = v$RD_7602_out0;
assign v$RD_6728_out0 = v$RD_7605_out0;
assign v$RD_6730_out0 = v$RD_7606_out0;
assign v$RD_6732_out0 = v$RD_7607_out0;
assign v$RD_6738_out0 = v$RD_7610_out0;
assign v$RD_6743_out0 = v$RD_7612_out0;
assign v$RD_6753_out0 = v$RD_7617_out0;
assign v$RD_6759_out0 = v$RD_7620_out0;
assign v$RD_6761_out0 = v$RD_7621_out0;
assign v$RD_6763_out0 = v$RD_7622_out0;
assign v$RD_6769_out0 = v$RD_7625_out0;
assign v$RD_6774_out0 = v$RD_7627_out0;
assign v$RD_6784_out0 = v$RD_7632_out0;
assign v$ADDER$IN_10995_out0 = v$_10783_out0;
assign v$NOTUSED_325_out0 = v$_3907_out0;
assign v$NOTUSED_326_out0 = v$_3908_out0;
assign v$ANDOUT_630_out0 = v$_1867_out0;
assign v$ANDOUT_632_out0 = v$_1869_out0;
assign v$_4483_out0 = v$MUX1_6_out0[1:0];
assign v$_4483_out1 = v$MUX1_6_out0[15:14];
assign v$_4484_out0 = v$MUX1_7_out0[1:0];
assign v$_4484_out1 = v$MUX1_7_out0[15:14];
assign v$_4591_out0 = { v$_3907_out1,v$C1_8815_out0 };
assign v$_4592_out0 = { v$_3908_out1,v$C1_8816_out0 };
assign v$_5846_out0 = v$A1_3174_out0[11:0];
assign v$_5846_out1 = v$A1_3174_out0[15:4];
assign v$_5847_out0 = v$A1_3175_out0[11:0];
assign v$_5847_out1 = v$A1_3175_out0[15:4];
assign v$COUT_10547_out0 = v$A1_3174_out1;
assign v$COUT_10548_out0 = v$A1_3175_out1;
assign v$RMN_13437_out0 = v$A1_3174_out0;
assign v$RMN_13438_out0 = v$A1_3175_out0;
assign v$OUT1_1972_out0 = v$_4591_out0;
assign v$OUT1_1973_out0 = v$_4592_out0;
assign v$NOTUSE_2399_out0 = v$_5846_out1;
assign v$NOTUSE_2400_out0 = v$_5847_out1;
assign v$_10910_out0 = v$ANDOUT_630_out0[0:0];
assign v$_10910_out1 = v$ANDOUT_630_out0[15:15];
assign v$_10911_out0 = v$ANDOUT_632_out0[0:0];
assign v$_10911_out1 = v$ANDOUT_632_out0[15:15];
assign v$UNUSED_11244_out0 = v$_4483_out0;
assign v$UNUSED_11245_out0 = v$_4484_out0;
assign v$_13482_out0 = { v$_4483_out1,v$C1_6793_out0 };
assign v$_13483_out0 = { v$_4484_out1,v$C1_6794_out0 };
assign v$MUX2_13656_out0 = v$G6_13258_out0 ? v$_5846_out0 : v$_3035_out0;
assign v$MUX2_13657_out0 = v$G6_13259_out0 ? v$_5847_out0 : v$_3036_out0;
assign v$CIN_2356_out0 = v$_10910_out1;
assign v$CIN_2371_out0 = v$_10911_out1;
assign v$MUX2_10841_out0 = v$LSR_13331_out0 ? v$_13482_out0 : v$MUX1_6_out0;
assign v$MUX2_10842_out0 = v$LSR_13332_out0 ? v$_13483_out0 : v$MUX1_7_out0;
assign v$EA_13516_out0 = v$MUX2_13656_out0;
assign v$EA_13517_out0 = v$MUX2_13657_out0;
assign v$MUX5_13670_out0 = v$0_3022_out0 ? v$OUT1_1972_out0 : v$IN_13668_out0;
assign v$MUX5_13671_out0 = v$0_3023_out0 ? v$OUT1_1973_out0 : v$IN_13669_out0;
assign v$_469_out0 = v$CIN_2356_out0[8:8];
assign v$_484_out0 = v$CIN_2371_out0[8:8];
assign v$_1774_out0 = v$CIN_2356_out0[6:6];
assign v$_1789_out0 = v$CIN_2371_out0[6:6];
assign v$IN_1964_out0 = v$MUX2_10841_out0;
assign v$IN_1965_out0 = v$MUX2_10842_out0;
assign v$_2156_out0 = v$CIN_2356_out0[3:3];
assign v$_2171_out0 = v$CIN_2371_out0[3:3];
assign v$RAMADDRMUX_2232_out0 = v$EA_13516_out0;
assign v$RAMADDRMUX_2233_out0 = v$EA_13517_out0;
assign v$_2503_out0 = v$CIN_2356_out0[0:0];
assign v$_2518_out0 = v$CIN_2371_out0[0:0];
assign v$_3052_out0 = v$CIN_2356_out0[9:9];
assign v$_3067_out0 = v$CIN_2371_out0[9:9];
assign v$_3086_out0 = v$CIN_2356_out0[2:2];
assign v$_3101_out0 = v$CIN_2371_out0[2:2];
assign v$_3140_out0 = v$CIN_2356_out0[7:7];
assign v$_3155_out0 = v$CIN_2371_out0[7:7];
assign v$_3824_out0 = v$CIN_2356_out0[1:1];
assign v$_3839_out0 = v$CIN_2371_out0[1:1];
assign v$_3862_out0 = v$CIN_2356_out0[10:10];
assign v$_3877_out0 = v$CIN_2371_out0[10:10];
assign v$_6801_out0 = v$CIN_2356_out0[11:11];
assign v$_6816_out0 = v$CIN_2371_out0[11:11];
assign v$_7645_out0 = v$CIN_2356_out0[12:12];
assign v$_7660_out0 = v$CIN_2371_out0[12:12];
assign v$_8700_out0 = v$CIN_2356_out0[13:13];
assign v$_8715_out0 = v$CIN_2371_out0[13:13];
assign v$_8770_out0 = v$CIN_2356_out0[14:14];
assign v$_8785_out0 = v$CIN_2371_out0[14:14];
assign v$_10720_out0 = v$CIN_2356_out0[5:5];
assign v$_10735_out0 = v$CIN_2371_out0[5:5];
assign v$IN1_10992_out0 = v$MUX5_13670_out0;
assign v$IN1_10993_out0 = v$MUX5_13671_out0;
assign v$_13449_out0 = v$CIN_2356_out0[4:4];
assign v$_13464_out0 = v$CIN_2371_out0[4:4];
assign v$RAMADDRMUX_92_out0 = v$RAMADDRMUX_2232_out0;
assign v$RAMADDRMUX_93_out0 = v$RAMADDRMUX_2233_out0;
assign v$_627_out0 = v$IN_1964_out0[1:0];
assign v$_627_out1 = v$IN_1964_out0[15:14];
assign v$_628_out0 = v$IN_1965_out0[1:0];
assign v$_628_out1 = v$IN_1965_out0[15:14];
assign v$RM_3370_out0 = v$_7645_out0;
assign v$RM_3371_out0 = v$_8770_out0;
assign v$RM_3372_out0 = v$_10720_out0;
assign v$RM_3373_out0 = v$_13449_out0;
assign v$RM_3374_out0 = v$_8700_out0;
assign v$RM_3375_out0 = v$_3052_out0;
assign v$RM_3376_out0 = v$_3862_out0;
assign v$RM_3377_out0 = v$_3824_out0;
assign v$RM_3378_out0 = v$_2156_out0;
assign v$RM_3379_out0 = v$_1774_out0;
assign v$RM_3380_out0 = v$_3140_out0;
assign v$RM_3381_out0 = v$_6801_out0;
assign v$RM_3382_out0 = v$_469_out0;
assign v$RM_3383_out0 = v$_3086_out0;
assign v$RM_3594_out0 = v$_7660_out0;
assign v$RM_3595_out0 = v$_8785_out0;
assign v$RM_3596_out0 = v$_10735_out0;
assign v$RM_3597_out0 = v$_13464_out0;
assign v$RM_3598_out0 = v$_8715_out0;
assign v$RM_3599_out0 = v$_3067_out0;
assign v$RM_3600_out0 = v$_3877_out0;
assign v$RM_3601_out0 = v$_3839_out0;
assign v$RM_3602_out0 = v$_2171_out0;
assign v$RM_3603_out0 = v$_1789_out0;
assign v$RM_3604_out0 = v$_3155_out0;
assign v$RM_3605_out0 = v$_6816_out0;
assign v$RM_3606_out0 = v$_484_out0;
assign v$RM_3607_out0 = v$_3101_out0;
assign v$_10823_out0 = v$IN_1964_out0[15:15];
assign v$_10824_out0 = v$IN_1965_out0[15:15];
assign v$RM_11343_out0 = v$_2503_out0;
assign v$RM_11807_out0 = v$_2518_out0;
assign v$_13550_out0 = v$IN1_10992_out0[1:0];
assign v$_13550_out1 = v$IN1_10992_out0[10:9];
assign v$_13551_out0 = v$IN1_10993_out0[1:0];
assign v$_13551_out1 = v$IN1_10993_out0[10:9];
assign v$NOTUSED_445_out0 = v$_13550_out0;
assign v$NOTUSED_446_out0 = v$_13551_out0;
assign v$NOTUSED_447_out0 = v$_627_out0;
assign v$NOTUSED_448_out0 = v$_628_out0;
assign v$G1_7758_out0 = ((v$RD_5903_out0 && !v$RM_11343_out0) || (!v$RD_5903_out0) && v$RM_11343_out0);
assign v$G1_8222_out0 = ((v$RD_6367_out0 && !v$RM_11807_out0) || (!v$RD_6367_out0) && v$RM_11807_out0);
assign v$_10354_out0 = { v$_627_out1,v$_10823_out0 };
assign v$_10355_out0 = { v$_628_out1,v$_10824_out0 };
assign v$RAMADDRMUX_10542_out0 = v$RAMADDRMUX_92_out0;
assign v$RAMADDRMUX_10543_out0 = v$RAMADDRMUX_93_out0;
assign v$RM_11333_out0 = v$RM_3370_out0;
assign v$RM_11335_out0 = v$RM_3371_out0;
assign v$RM_11337_out0 = v$RM_3372_out0;
assign v$RM_11339_out0 = v$RM_3373_out0;
assign v$RM_11341_out0 = v$RM_3374_out0;
assign v$RM_11345_out0 = v$RM_3375_out0;
assign v$RM_11347_out0 = v$RM_3376_out0;
assign v$RM_11349_out0 = v$RM_3377_out0;
assign v$RM_11351_out0 = v$RM_3378_out0;
assign v$RM_11353_out0 = v$RM_3379_out0;
assign v$RM_11355_out0 = v$RM_3380_out0;
assign v$RM_11357_out0 = v$RM_3381_out0;
assign v$RM_11359_out0 = v$RM_3382_out0;
assign v$RM_11361_out0 = v$RM_3383_out0;
assign v$RM_11797_out0 = v$RM_3594_out0;
assign v$RM_11799_out0 = v$RM_3595_out0;
assign v$RM_11801_out0 = v$RM_3596_out0;
assign v$RM_11803_out0 = v$RM_3597_out0;
assign v$RM_11805_out0 = v$RM_3598_out0;
assign v$RM_11809_out0 = v$RM_3599_out0;
assign v$RM_11811_out0 = v$RM_3600_out0;
assign v$RM_11813_out0 = v$RM_3601_out0;
assign v$RM_11815_out0 = v$RM_3602_out0;
assign v$RM_11817_out0 = v$RM_3603_out0;
assign v$RM_11819_out0 = v$RM_3604_out0;
assign v$RM_11821_out0 = v$RM_3605_out0;
assign v$RM_11823_out0 = v$RM_3606_out0;
assign v$RM_11825_out0 = v$RM_3607_out0;
assign v$G2_12294_out0 = v$RD_5903_out0 && v$RM_11343_out0;
assign v$G2_12758_out0 = v$RD_6367_out0 && v$RM_11807_out0;
assign v$_13761_out0 = { v$_13550_out1,v$C1_3205_out0 };
assign v$_13762_out0 = { v$_13551_out1,v$C1_3206_out0 };
assign v$_1172_out0 = { v$_10354_out0,v$_10823_out0 };
assign v$_1173_out0 = { v$_10355_out0,v$_10824_out0 };
assign v$OUT1_3853_out0 = v$_13761_out0;
assign v$OUT1_3854_out0 = v$_13762_out0;
assign v$CARRY_4903_out0 = v$G2_12294_out0;
assign v$CARRY_5367_out0 = v$G2_12758_out0;
assign v$G1_7748_out0 = ((v$RD_5893_out0 && !v$RM_11333_out0) || (!v$RD_5893_out0) && v$RM_11333_out0);
assign v$G1_7750_out0 = ((v$RD_5895_out0 && !v$RM_11335_out0) || (!v$RD_5895_out0) && v$RM_11335_out0);
assign v$G1_7752_out0 = ((v$RD_5897_out0 && !v$RM_11337_out0) || (!v$RD_5897_out0) && v$RM_11337_out0);
assign v$G1_7754_out0 = ((v$RD_5899_out0 && !v$RM_11339_out0) || (!v$RD_5899_out0) && v$RM_11339_out0);
assign v$G1_7756_out0 = ((v$RD_5901_out0 && !v$RM_11341_out0) || (!v$RD_5901_out0) && v$RM_11341_out0);
assign v$G1_7760_out0 = ((v$RD_5905_out0 && !v$RM_11345_out0) || (!v$RD_5905_out0) && v$RM_11345_out0);
assign v$G1_7762_out0 = ((v$RD_5907_out0 && !v$RM_11347_out0) || (!v$RD_5907_out0) && v$RM_11347_out0);
assign v$G1_7764_out0 = ((v$RD_5909_out0 && !v$RM_11349_out0) || (!v$RD_5909_out0) && v$RM_11349_out0);
assign v$G1_7766_out0 = ((v$RD_5911_out0 && !v$RM_11351_out0) || (!v$RD_5911_out0) && v$RM_11351_out0);
assign v$G1_7768_out0 = ((v$RD_5913_out0 && !v$RM_11353_out0) || (!v$RD_5913_out0) && v$RM_11353_out0);
assign v$G1_7770_out0 = ((v$RD_5915_out0 && !v$RM_11355_out0) || (!v$RD_5915_out0) && v$RM_11355_out0);
assign v$G1_7772_out0 = ((v$RD_5917_out0 && !v$RM_11357_out0) || (!v$RD_5917_out0) && v$RM_11357_out0);
assign v$G1_7774_out0 = ((v$RD_5919_out0 && !v$RM_11359_out0) || (!v$RD_5919_out0) && v$RM_11359_out0);
assign v$G1_7776_out0 = ((v$RD_5921_out0 && !v$RM_11361_out0) || (!v$RD_5921_out0) && v$RM_11361_out0);
assign v$G1_8212_out0 = ((v$RD_6357_out0 && !v$RM_11797_out0) || (!v$RD_6357_out0) && v$RM_11797_out0);
assign v$G1_8214_out0 = ((v$RD_6359_out0 && !v$RM_11799_out0) || (!v$RD_6359_out0) && v$RM_11799_out0);
assign v$G1_8216_out0 = ((v$RD_6361_out0 && !v$RM_11801_out0) || (!v$RD_6361_out0) && v$RM_11801_out0);
assign v$G1_8218_out0 = ((v$RD_6363_out0 && !v$RM_11803_out0) || (!v$RD_6363_out0) && v$RM_11803_out0);
assign v$G1_8220_out0 = ((v$RD_6365_out0 && !v$RM_11805_out0) || (!v$RD_6365_out0) && v$RM_11805_out0);
assign v$G1_8224_out0 = ((v$RD_6369_out0 && !v$RM_11809_out0) || (!v$RD_6369_out0) && v$RM_11809_out0);
assign v$G1_8226_out0 = ((v$RD_6371_out0 && !v$RM_11811_out0) || (!v$RD_6371_out0) && v$RM_11811_out0);
assign v$G1_8228_out0 = ((v$RD_6373_out0 && !v$RM_11813_out0) || (!v$RD_6373_out0) && v$RM_11813_out0);
assign v$G1_8230_out0 = ((v$RD_6375_out0 && !v$RM_11815_out0) || (!v$RD_6375_out0) && v$RM_11815_out0);
assign v$G1_8232_out0 = ((v$RD_6377_out0 && !v$RM_11817_out0) || (!v$RD_6377_out0) && v$RM_11817_out0);
assign v$G1_8234_out0 = ((v$RD_6379_out0 && !v$RM_11819_out0) || (!v$RD_6379_out0) && v$RM_11819_out0);
assign v$G1_8236_out0 = ((v$RD_6381_out0 && !v$RM_11821_out0) || (!v$RD_6381_out0) && v$RM_11821_out0);
assign v$G1_8238_out0 = ((v$RD_6383_out0 && !v$RM_11823_out0) || (!v$RD_6383_out0) && v$RM_11823_out0);
assign v$G1_8240_out0 = ((v$RD_6385_out0 && !v$RM_11825_out0) || (!v$RD_6385_out0) && v$RM_11825_out0);
assign v$RAM$ADDRESS$MUX_8803_out0 = v$RAMADDRMUX_10542_out0;
assign v$RAM$ADDRESS$MUX_8804_out0 = v$RAMADDRMUX_10543_out0;
assign v$S_8904_out0 = v$G1_7758_out0;
assign v$S_9368_out0 = v$G1_8222_out0;
assign v$G2_12284_out0 = v$RD_5893_out0 && v$RM_11333_out0;
assign v$G2_12286_out0 = v$RD_5895_out0 && v$RM_11335_out0;
assign v$G2_12288_out0 = v$RD_5897_out0 && v$RM_11337_out0;
assign v$G2_12290_out0 = v$RD_5899_out0 && v$RM_11339_out0;
assign v$G2_12292_out0 = v$RD_5901_out0 && v$RM_11341_out0;
assign v$G2_12296_out0 = v$RD_5905_out0 && v$RM_11345_out0;
assign v$G2_12298_out0 = v$RD_5907_out0 && v$RM_11347_out0;
assign v$G2_12300_out0 = v$RD_5909_out0 && v$RM_11349_out0;
assign v$G2_12302_out0 = v$RD_5911_out0 && v$RM_11351_out0;
assign v$G2_12304_out0 = v$RD_5913_out0 && v$RM_11353_out0;
assign v$G2_12306_out0 = v$RD_5915_out0 && v$RM_11355_out0;
assign v$G2_12308_out0 = v$RD_5917_out0 && v$RM_11357_out0;
assign v$G2_12310_out0 = v$RD_5919_out0 && v$RM_11359_out0;
assign v$G2_12312_out0 = v$RD_5921_out0 && v$RM_11361_out0;
assign v$G2_12748_out0 = v$RD_6357_out0 && v$RM_11797_out0;
assign v$G2_12750_out0 = v$RD_6359_out0 && v$RM_11799_out0;
assign v$G2_12752_out0 = v$RD_6361_out0 && v$RM_11801_out0;
assign v$G2_12754_out0 = v$RD_6363_out0 && v$RM_11803_out0;
assign v$G2_12756_out0 = v$RD_6365_out0 && v$RM_11805_out0;
assign v$G2_12760_out0 = v$RD_6369_out0 && v$RM_11809_out0;
assign v$G2_12762_out0 = v$RD_6371_out0 && v$RM_11811_out0;
assign v$G2_12764_out0 = v$RD_6373_out0 && v$RM_11813_out0;
assign v$G2_12766_out0 = v$RD_6375_out0 && v$RM_11815_out0;
assign v$G2_12768_out0 = v$RD_6377_out0 && v$RM_11817_out0;
assign v$G2_12770_out0 = v$RD_6379_out0 && v$RM_11819_out0;
assign v$G2_12772_out0 = v$RD_6381_out0 && v$RM_11821_out0;
assign v$G2_12774_out0 = v$RD_6383_out0 && v$RM_11823_out0;
assign v$G2_12776_out0 = v$RD_6385_out0 && v$RM_11825_out0;
assign v$RAM$ADDRES$MUX_13649_out0 = v$RAMADDRMUX_10542_out0;
assign v$RAM$ADDRES$MUX_13650_out0 = v$RAMADDRMUX_10543_out0;
assign v$MUX4_552_out0 = v$1_3817_out0 ? v$OUT1_3853_out0 : v$MUX5_13670_out0;
assign v$MUX4_553_out0 = v$1_3818_out0 ? v$OUT1_3854_out0 : v$MUX5_13671_out0;
assign v$ADRESS1_1906_out0 = v$RAM$ADDRES$MUX_13649_out0;
assign v$S_4666_out0 = v$S_8904_out0;
assign v$S_4681_out0 = v$S_9368_out0;
assign v$CARRY_4893_out0 = v$G2_12284_out0;
assign v$CARRY_4895_out0 = v$G2_12286_out0;
assign v$CARRY_4897_out0 = v$G2_12288_out0;
assign v$CARRY_4899_out0 = v$G2_12290_out0;
assign v$CARRY_4901_out0 = v$G2_12292_out0;
assign v$CARRY_4905_out0 = v$G2_12296_out0;
assign v$CARRY_4907_out0 = v$G2_12298_out0;
assign v$CARRY_4909_out0 = v$G2_12300_out0;
assign v$CARRY_4911_out0 = v$G2_12302_out0;
assign v$CARRY_4913_out0 = v$G2_12304_out0;
assign v$CARRY_4915_out0 = v$G2_12306_out0;
assign v$CARRY_4917_out0 = v$G2_12308_out0;
assign v$CARRY_4919_out0 = v$G2_12310_out0;
assign v$CARRY_4921_out0 = v$G2_12312_out0;
assign v$CARRY_5357_out0 = v$G2_12748_out0;
assign v$CARRY_5359_out0 = v$G2_12750_out0;
assign v$CARRY_5361_out0 = v$G2_12752_out0;
assign v$CARRY_5363_out0 = v$G2_12754_out0;
assign v$CARRY_5365_out0 = v$G2_12756_out0;
assign v$CARRY_5369_out0 = v$G2_12760_out0;
assign v$CARRY_5371_out0 = v$G2_12762_out0;
assign v$CARRY_5373_out0 = v$G2_12764_out0;
assign v$CARRY_5375_out0 = v$G2_12766_out0;
assign v$CARRY_5377_out0 = v$G2_12768_out0;
assign v$CARRY_5379_out0 = v$G2_12770_out0;
assign v$CARRY_5381_out0 = v$G2_12772_out0;
assign v$CARRY_5383_out0 = v$G2_12774_out0;
assign v$CARRY_5385_out0 = v$G2_12776_out0;
assign v$RAMADDRMUX_7066_out0 = v$RAM$ADDRESS$MUX_8803_out0;
assign v$RAMADDRMUX_7067_out0 = v$RAM$ADDRESS$MUX_8804_out0;
assign v$OUT_8852_out0 = v$_1172_out0;
assign v$OUT_8853_out0 = v$_1173_out0;
assign v$S_8894_out0 = v$G1_7748_out0;
assign v$S_8896_out0 = v$G1_7750_out0;
assign v$S_8898_out0 = v$G1_7752_out0;
assign v$S_8900_out0 = v$G1_7754_out0;
assign v$S_8902_out0 = v$G1_7756_out0;
assign v$S_8906_out0 = v$G1_7760_out0;
assign v$S_8908_out0 = v$G1_7762_out0;
assign v$S_8910_out0 = v$G1_7764_out0;
assign v$S_8912_out0 = v$G1_7766_out0;
assign v$S_8914_out0 = v$G1_7768_out0;
assign v$S_8916_out0 = v$G1_7770_out0;
assign v$S_8918_out0 = v$G1_7772_out0;
assign v$S_8920_out0 = v$G1_7774_out0;
assign v$S_8922_out0 = v$G1_7776_out0;
assign v$S_9358_out0 = v$G1_8212_out0;
assign v$S_9360_out0 = v$G1_8214_out0;
assign v$S_9362_out0 = v$G1_8216_out0;
assign v$S_9364_out0 = v$G1_8218_out0;
assign v$S_9366_out0 = v$G1_8220_out0;
assign v$S_9370_out0 = v$G1_8224_out0;
assign v$S_9372_out0 = v$G1_8226_out0;
assign v$S_9374_out0 = v$G1_8228_out0;
assign v$S_9376_out0 = v$G1_8230_out0;
assign v$S_9378_out0 = v$G1_8232_out0;
assign v$S_9380_out0 = v$G1_8234_out0;
assign v$S_9382_out0 = v$G1_8236_out0;
assign v$S_9384_out0 = v$G1_8238_out0;
assign v$S_9386_out0 = v$G1_8240_out0;
assign v$CIN_9830_out0 = v$CARRY_4903_out0;
assign v$CIN_10054_out0 = v$CARRY_5367_out0;
assign v$ADRESS0_11217_out0 = v$RAM$ADDRES$MUX_13650_out0;
assign v$_2437_out0 = v$RAMADDRMUX_7066_out0[3:0];
assign v$_2437_out1 = v$RAMADDRMUX_7066_out0[11:8];
assign v$_2438_out0 = v$RAMADDRMUX_7067_out0[3:0];
assign v$_2438_out1 = v$RAMADDRMUX_7067_out0[11:8];
assign v$IN1_2848_out0 = v$MUX4_552_out0;
assign v$IN1_2849_out0 = v$MUX4_553_out0;
assign v$ADDRESS1_2854_out0 = v$ADRESS1_1906_out0;
assign v$MUX3_3133_out0 = v$ASR_13713_out0 ? v$OUT_8852_out0 : v$MUX2_10841_out0;
assign v$MUX3_3134_out0 = v$ASR_13714_out0 ? v$OUT_8853_out0 : v$MUX2_10842_out0;
assign v$_3223_out0 = { v$_10910_out0,v$S_4666_out0 };
assign v$_3224_out0 = { v$_10911_out0,v$S_4681_out0 };
assign v$EQ11_4465_out0 = v$RAMADDRMUX_7066_out0 == 12'h800;
assign v$EQ11_4466_out0 = v$RAMADDRMUX_7067_out0 == 12'h800;
assign v$RD_5910_out0 = v$CIN_9830_out0;
assign v$RD_6374_out0 = v$CIN_10054_out0;
assign v$ADDRESS0_10982_out0 = v$ADRESS0_11217_out0;
assign v$RM_11334_out0 = v$S_8894_out0;
assign v$RM_11336_out0 = v$S_8896_out0;
assign v$RM_11338_out0 = v$S_8898_out0;
assign v$RM_11340_out0 = v$S_8900_out0;
assign v$RM_11342_out0 = v$S_8902_out0;
assign v$RM_11346_out0 = v$S_8906_out0;
assign v$RM_11348_out0 = v$S_8908_out0;
assign v$RM_11350_out0 = v$S_8910_out0;
assign v$RM_11352_out0 = v$S_8912_out0;
assign v$RM_11354_out0 = v$S_8914_out0;
assign v$RM_11356_out0 = v$S_8916_out0;
assign v$RM_11358_out0 = v$S_8918_out0;
assign v$RM_11360_out0 = v$S_8920_out0;
assign v$RM_11362_out0 = v$S_8922_out0;
assign v$RM_11798_out0 = v$S_9358_out0;
assign v$RM_11800_out0 = v$S_9360_out0;
assign v$RM_11802_out0 = v$S_9362_out0;
assign v$RM_11804_out0 = v$S_9364_out0;
assign v$RM_11806_out0 = v$S_9366_out0;
assign v$RM_11810_out0 = v$S_9370_out0;
assign v$RM_11812_out0 = v$S_9372_out0;
assign v$RM_11814_out0 = v$S_9374_out0;
assign v$RM_11816_out0 = v$S_9376_out0;
assign v$RM_11818_out0 = v$S_9378_out0;
assign v$RM_11820_out0 = v$S_9380_out0;
assign v$RM_11822_out0 = v$S_9382_out0;
assign v$RM_11824_out0 = v$S_9384_out0;
assign v$RM_11826_out0 = v$S_9386_out0;
assign v$_4703_out0 = v$IN1_2848_out0[3:0];
assign v$_4703_out1 = v$IN1_2848_out0[10:7];
assign v$_4704_out0 = v$IN1_2849_out0[3:0];
assign v$_4704_out1 = v$IN1_2849_out0[10:7];
assign v$_4816_out0 = v$MUX3_3133_out0[1:0];
assign v$_4816_out1 = v$MUX3_3133_out0[15:14];
assign v$_4817_out0 = v$MUX3_3134_out0[1:0];
assign v$_4817_out1 = v$MUX3_3134_out0[15:14];
assign v$MUX1_7097_out0 = v$MUX$ENABLE_2349_out0 ? v$ADDRESS0_10982_out0 : v$ADDRESS1_2854_out0;
assign v$G1_7765_out0 = ((v$RD_5910_out0 && !v$RM_11350_out0) || (!v$RD_5910_out0) && v$RM_11350_out0);
assign v$G1_8229_out0 = ((v$RD_6374_out0 && !v$RM_11814_out0) || (!v$RD_6374_out0) && v$RM_11814_out0);
assign v$G2_12301_out0 = v$RD_5910_out0 && v$RM_11350_out0;
assign v$G2_12765_out0 = v$RD_6374_out0 && v$RM_11814_out0;
assign v$_13317_out0 = v$_2437_out1[3:0];
assign v$_13317_out1 = v$_2437_out1[7:4];
assign v$_13318_out0 = v$_2438_out1[3:0];
assign v$_13318_out1 = v$_2438_out1[7:4];
assign v$RAM$ADD$BYTE0_13382_out0 = v$_2437_out0;
assign v$RAM$ADD$BYTE0_13383_out0 = v$_2438_out0;
assign v$G22_13707_out0 = v$EQ11_4465_out0 && v$UART_11128_out0;
assign v$G22_13708_out0 = v$EQ11_4466_out0 && v$UART_11129_out0;
assign v$_1209_out0 = { v$_4816_out1,v$_4816_out0 };
assign v$_1210_out0 = { v$_4817_out1,v$_4817_out0 };
assign v$EQ1_2675_out0 = v$_13317_out0 == 4'h1;
assign v$EQ1_2676_out0 = v$_13318_out0 == 4'h1;
assign v$_2971_out0 = { v$_4703_out1,v$C1_10305_out0 };
assign v$_2972_out0 = { v$_4704_out1,v$C1_10306_out0 };
assign v$ADDRESS_4662_out0 = v$MUX1_7097_out0;
assign v$EQ9_4842_out0 = v$RAM$ADD$BYTE0_13382_out0 == 4'h2;
assign v$EQ9_4843_out0 = v$RAM$ADD$BYTE0_13383_out0 == 4'h2;
assign v$CARRY_4910_out0 = v$G2_12301_out0;
assign v$CARRY_5374_out0 = v$G2_12765_out0;
assign v$S_8911_out0 = v$G1_7765_out0;
assign v$S_9375_out0 = v$G1_8229_out0;
assign v$G23_10439_out0 = v$G22_13707_out0 && v$LOAD_3949_out0;
assign v$G23_10440_out0 = v$G22_13708_out0 && v$LOAD_3950_out0;
assign v$EQ01_10510_out0 = v$RAM$ADD$BYTE0_13382_out0 == 4'h1;
assign v$EQ01_10511_out0 = v$RAM$ADD$BYTE0_13383_out0 == 4'h1;
assign v$NOTUSED_10540_out0 = v$_4703_out0;
assign v$NOTUSED_10541_out0 = v$_4704_out0;
assign v$EQ8_10804_out0 = v$_13317_out1 == 4'h8;
assign v$EQ8_10805_out0 = v$_13318_out1 == 4'h8;
assign v$S_1241_out0 = v$S_8911_out0;
assign v$S_1465_out0 = v$S_9375_out0;
assign v$OUT1_1873_out0 = v$_2971_out0;
assign v$OUT1_1874_out0 = v$_2972_out0;
assign v$BYTE1$comp1_2443_out0 = v$EQ1_2675_out0;
assign v$BYTE1$comp1_2444_out0 = v$EQ1_2676_out0;
assign v$STAT$INSTRUCTION_2855_out0 = v$G23_10439_out0;
assign v$STAT$INSTRUCTION_2856_out0 = v$G23_10440_out0;
assign v$G1_4017_out0 = v$CARRY_4910_out0 || v$CARRY_4909_out0;
assign v$G1_4241_out0 = v$CARRY_5374_out0 || v$CARRY_5373_out0;
assign v$BYTE2$COMP8_7695_out0 = v$EQ8_10804_out0;
assign v$BYTE2$COMP8_7696_out0 = v$EQ8_10805_out0;
assign v$ADRESS_8683_out0 = v$ADDRESS_4662_out0;
assign v$MUX4_10524_out0 = v$ROR_3286_out0 ? v$_1209_out0 : v$MUX3_3133_out0;
assign v$MUX4_10525_out0 = v$ROR_3287_out0 ? v$_1210_out0 : v$MUX3_3134_out0;
assign v$COUT_709_out0 = v$G1_4017_out0;
assign v$COUT_933_out0 = v$G1_4241_out0;
assign v$MUX5_1185_out0 = v$EN_10474_out0 ? v$MUX4_10524_out0 : v$IN_8838_out0;
assign v$MUX5_1186_out0 = v$EN_10475_out0 ? v$MUX4_10525_out0 : v$IN_8839_out0;
assign v$STAT$INSTRUCTION_2434_out0 = v$STAT$INSTRUCTION_2855_out0;
assign v$STAT$INSTRUCTION_2435_out0 = v$STAT$INSTRUCTION_2856_out0;
assign v$G2_3245_out0 = v$EQ01_10510_out0 && v$BYTE2$COMP8_7695_out0;
assign v$G2_3246_out0 = v$EQ01_10511_out0 && v$BYTE2$COMP8_7696_out0;
assign v$BYTE$COMP1_3262_out0 = v$BYTE1$comp1_2443_out0;
assign v$BYTE$COMP1_3263_out0 = v$BYTE1$comp1_2444_out0;
assign v$G20_11147_out0 = v$BYTE2$COMP8_7695_out0 && v$EQ9_4842_out0;
assign v$G20_11148_out0 = v$BYTE2$COMP8_7696_out0 && v$EQ9_4843_out0;
assign v$MUX3_13312_out0 = v$2_1763_out0 ? v$OUT1_1873_out0 : v$MUX4_552_out0;
assign v$MUX3_13313_out0 = v$2_1764_out0 ? v$OUT1_1874_out0 : v$MUX4_553_out0;
assign v$MUX3_13335_out0 = v$BYTE1$comp1_2443_out0 ? v$_9791_out0 : v$_7081_out0;
assign v$MUX3_13336_out0 = v$BYTE1$comp1_2444_out0 ? v$_9792_out0 : v$_7082_out0;
assign v$BYTE$COMP1_9796_out0 = v$BYTE$COMP1_3262_out0;
assign v$BYTE$COMP1_9797_out0 = v$BYTE$COMP1_3263_out0;
assign v$CIN_9836_out0 = v$COUT_709_out0;
assign v$CIN_10060_out0 = v$COUT_933_out0;
assign v$STAT$INSTRUCTION_10272_out0 = v$STAT$INSTRUCTION_2434_out0;
assign v$STAT$INSTRUCTION_10273_out0 = v$STAT$INSTRUCTION_2435_out0;
assign v$G14_10407_out0 = v$G2_3245_out0 && v$UART_11128_out0;
assign v$G14_10408_out0 = v$G2_3246_out0 && v$UART_11129_out0;
assign v$G18_11204_out0 = v$G20_11147_out0 && v$UART_11128_out0;
assign v$G18_11205_out0 = v$G20_11148_out0 && v$UART_11129_out0;
assign v$OUT_12236_out0 = v$MUX5_1185_out0;
assign v$OUT_12237_out0 = v$MUX5_1186_out0;
assign v$IN1_13711_out0 = v$MUX3_13312_out0;
assign v$IN1_13712_out0 = v$MUX3_13313_out0;
assign v$byte$comp$10_2318_out0 = v$BYTE$COMP1_9797_out0;
assign v$byte$comp$11_2645_out0 = v$BYTE$COMP1_9796_out0;
assign v$IN_2664_out0 = v$OUT_12236_out0;
assign v$IN_2665_out0 = v$OUT_12237_out0;
assign v$_2680_out0 = v$IN1_13711_out0[7:0];
assign v$_2680_out1 = v$IN1_13711_out0[10:3];
assign v$_2681_out0 = v$IN1_13712_out0[7:0];
assign v$_2681_out1 = v$IN1_13712_out0[10:3];
assign v$G19_4663_out0 = v$G18_11204_out0 && v$STORE_221_out0;
assign v$G19_4664_out0 = v$G18_11205_out0 && v$STORE_222_out0;
assign v$RD_5922_out0 = v$CIN_9836_out0;
assign v$RD_6386_out0 = v$CIN_10060_out0;
assign v$G16_13388_out0 = v$G14_10407_out0 && v$LOAD_3949_out0;
assign v$G16_13389_out0 = v$G14_10408_out0 && v$LOAD_3950_out0;
assign v$NOTUSED_683_out0 = v$_2680_out0;
assign v$NOTUSED_684_out0 = v$_2681_out0;
assign v$BYTE$COMP$11_1163_out0 = v$byte$comp$11_2645_out0;
assign v$_2411_out0 = v$IN_2664_out0[11:0];
assign v$_2411_out1 = v$IN_2664_out0[15:4];
assign v$_2412_out0 = v$IN_2665_out0[11:0];
assign v$_2412_out1 = v$IN_2665_out0[15:4];
assign v$G21_2885_out0 = v$G19_4663_out0 && v$EXEC1_3038_out0;
assign v$G21_2886_out0 = v$G19_4664_out0 && v$EXEC1_3039_out0;
assign v$G1_7777_out0 = ((v$RD_5922_out0 && !v$RM_11362_out0) || (!v$RD_5922_out0) && v$RM_11362_out0);
assign v$G1_8241_out0 = ((v$RD_6386_out0 && !v$RM_11826_out0) || (!v$RD_6386_out0) && v$RM_11826_out0);
assign v$RX$INSTRUCTION_11170_out0 = v$G16_13388_out0;
assign v$RX$INSTRUCTION_11171_out0 = v$G16_13389_out0;
assign v$G2_12313_out0 = v$RD_5922_out0 && v$RM_11362_out0;
assign v$G2_12777_out0 = v$RD_6386_out0 && v$RM_11826_out0;
assign v$_13484_out0 = { v$_2680_out1,v$C1_10266_out0 };
assign v$_13485_out0 = { v$_2681_out1,v$C1_10267_out0 };
assign v$IN_13548_out0 = v$IN_2664_out0;
assign v$IN_13549_out0 = v$IN_2665_out0;
assign v$BYTE$COMP$10_13611_out0 = v$byte$comp$10_2318_out0;
assign v$TX$INSTRUCTION_62_out0 = v$G21_2885_out0;
assign v$TX$INSTRUCTION_63_out0 = v$G21_2886_out0;
assign v$RX$INSTRUCTION_94_out0 = v$RX$INSTRUCTION_11170_out0;
assign v$RX$INSTRUCTION_95_out0 = v$RX$INSTRUCTION_11171_out0;
assign v$NOTUSED1_1897_out0 = v$_2411_out1;
assign v$NOTUSED1_1898_out0 = v$_2412_out1;
assign v$_2678_out0 = { v$C1_6919_out0,v$_2411_out0 };
assign v$_2679_out0 = { v$C1_6920_out0,v$_2412_out0 };
assign v$OUT1_3294_out0 = v$_13484_out0;
assign v$OUT1_3295_out0 = v$_13485_out0;
assign v$CARRY_4922_out0 = v$G2_12313_out0;
assign v$CARRY_5386_out0 = v$G2_12777_out0;
assign v$S_8923_out0 = v$G1_7777_out0;
assign v$S_9387_out0 = v$G1_8241_out0;
assign v$MUX1_11141_out0 = v$RX$INSTRUCTION_11170_out0 ? v$MUX3_13335_out0 : v$RAM$OUT_11214_out0;
assign v$MUX1_11142_out0 = v$RX$INSTRUCTION_11171_out0 ? v$MUX3_13336_out0 : v$RAM$OUT_11215_out0;
assign v$S_1247_out0 = v$S_8923_out0;
assign v$S_1471_out0 = v$S_9387_out0;
assign v$RX$INSTRUCTION_3258_out0 = v$RX$INSTRUCTION_94_out0;
assign v$RX$INSTRUCTION_3259_out0 = v$RX$INSTRUCTION_95_out0;
assign v$G1_4023_out0 = v$CARRY_4922_out0 || v$CARRY_4921_out0;
assign v$G1_4247_out0 = v$CARRY_5386_out0 || v$CARRY_5385_out0;
assign v$MUX1_4844_out0 = v$LSL_3047_out0 ? v$_2678_out0 : v$IN_13548_out0;
assign v$MUX1_4845_out0 = v$LSL_3048_out0 ? v$_2679_out0 : v$IN_13549_out0;
assign v$TX$INSTRUCTION_7012_out0 = v$TX$INSTRUCTION_62_out0;
assign v$TX$INSTRUCTION_7013_out0 = v$TX$INSTRUCTION_63_out0;
assign v$MUX1_7143_out0 = v$3_13619_out0 ? v$OUT1_3294_out0 : v$MUX3_13312_out0;
assign v$MUX1_7144_out0 = v$3_13620_out0 ? v$OUT1_3295_out0 : v$MUX3_13313_out0;
assign v$REGISTER$INPUT_13270_out0 = v$MUX1_11141_out0;
assign v$REGISTER$INPUT_13271_out0 = v$MUX1_11142_out0;
assign v$COUT_715_out0 = v$G1_4023_out0;
assign v$COUT_939_out0 = v$G1_4247_out0;
assign v$RX$INSTRUCTION_2343_out0 = v$RX$INSTRUCTION_3258_out0;
assign v$RX$INSTRUCTION_2344_out0 = v$RX$INSTRUCTION_3259_out0;
assign v$shifted1_2666_out0 = v$MUX1_7143_out0;
assign v$shifted1_2667_out0 = v$MUX1_7144_out0;
assign v$REGISTE$IN_4490_out0 = v$REGISTER$INPUT_13270_out0;
assign v$REGISTE$IN_4491_out0 = v$REGISTER$INPUT_13271_out0;
assign v$_4585_out0 = v$MUX1_4844_out0[3:0];
assign v$_4585_out1 = v$MUX1_4844_out0[15:12];
assign v$_4586_out0 = v$MUX1_4845_out0[3:0];
assign v$_4586_out1 = v$MUX1_4845_out0[15:12];
assign v$_4783_out0 = { v$S_1241_out0,v$S_1247_out0 };
assign v$_4798_out0 = { v$S_1465_out0,v$S_1471_out0 };
assign v$TX$INSTRUCTION_13659_out0 = v$TX$INSTRUCTION_7012_out0;
assign v$TX$INSTRUCTION_13660_out0 = v$TX$INSTRUCTION_7013_out0;
assign v$RX$INST1_12_out0 = v$RX$INSTRUCTION_2343_out0;
assign v$RX$INST0_2970_out0 = v$RX$INSTRUCTION_2344_out0;
assign v$RAMDOUT_3031_out0 = v$REGISTE$IN_4490_out0;
assign v$RAMDOUT_3032_out0 = v$REGISTE$IN_4491_out0;
assign v$_4660_out0 = { v$_4585_out1,v$C1_6919_out0 };
assign v$_4661_out0 = { v$_4586_out1,v$C1_6920_out0 };
assign v$NOTUSED_9800_out0 = v$_4585_out0;
assign v$NOTUSED_9801_out0 = v$_4586_out0;
assign v$CIN_9831_out0 = v$COUT_715_out0;
assign v$CIN_10055_out0 = v$COUT_939_out0;
assign v$TX$INST_10827_out0 = v$TX$INSTRUCTION_13659_out0;
assign v$TX$INST_10828_out0 = v$TX$INSTRUCTION_13660_out0;
assign v$REGISTER$INPUT_13621_out0 = v$REGISTE$IN_4490_out0;
assign v$REGISTER$INPUT_13622_out0 = v$REGISTE$IN_4491_out0;
assign v$SHIFTED$SIG_13632_out0 = v$shifted1_2666_out0;
assign v$SHIFTED$SIG_13633_out0 = v$shifted1_2667_out0;
assign v$RAMDOUT_23_out0 = v$RAMDOUT_3031_out0;
assign v$RAMDOUT_24_out0 = v$RAMDOUT_3032_out0;
assign v$REGISTER$INUP16_384_out0 = v$REGISTER$INPUT_13621_out0;
assign v$TX$INSTRUCTION1_1169_out0 = v$TX$INST_10827_out0;
assign v$TX$INSTRUCTION0_1762_out0 = v$TX$INST_10828_out0;
assign v$G1_2354_out0 = v$RX$INST1_12_out0 || v$RX$INST0_2970_out0;
assign v$RD_5912_out0 = v$CIN_9831_out0;
assign v$RD_6376_out0 = v$CIN_10055_out0;
assign v$SHIFTED$SIG_10802_out0 = v$SHIFTED$SIG_13632_out0;
assign v$SHIFTED$SIG_10803_out0 = v$SHIFTED$SIG_13633_out0;
assign v$REGISTER$INUP0_12240_out0 = v$REGISTER$INPUT_13622_out0;
assign v$MUX2_13319_out0 = v$LSR_418_out0 ? v$_4660_out0 : v$MUX1_4844_out0;
assign v$MUX2_13320_out0 = v$LSR_419_out0 ? v$_4661_out0 : v$MUX1_4845_out0;
assign v$MUX2_188_out0 = v$SHIFT$WHICH$OP_4459_out0 ? v$RD$SIG11_7132_out0 : v$SHIFTED$SIG_10802_out0;
assign v$MUX2_189_out0 = v$SHIFT$WHICH$OP_4460_out0 ? v$RD$SIG11_7133_out0 : v$SHIFTED$SIG_10803_out0;
assign v$TX$INSTUCTION0_228_out0 = v$TX$INSTRUCTION0_1762_out0;
assign v$RX$INST_2334_out0 = v$G1_2354_out0;
assign v$IN_2350_out0 = v$MUX2_13319_out0;
assign v$IN_2351_out0 = v$MUX2_13320_out0;
assign v$RAMDOUT_2414_out0 = v$RAMDOUT_23_out0;
assign v$RAMDOUT_2415_out0 = v$RAMDOUT_24_out0;
assign v$TX$INSTUCTION1_4859_out0 = v$TX$INSTRUCTION1_1169_out0;
assign v$MUX1_7702_out0 = v$SHIFT$WHICH$OP_4459_out0 ? v$SHIFTED$SIG_10802_out0 : v$OP2$SIG11_4827_out0;
assign v$MUX1_7703_out0 = v$SHIFT$WHICH$OP_4460_out0 ? v$SHIFTED$SIG_10803_out0 : v$OP2$SIG11_4828_out0;
assign v$G1_7767_out0 = ((v$RD_5912_out0 && !v$RM_11352_out0) || (!v$RD_5912_out0) && v$RM_11352_out0);
assign v$G1_8231_out0 = ((v$RD_6376_out0 && !v$RM_11816_out0) || (!v$RD_6376_out0) && v$RM_11816_out0);
assign v$G2_12303_out0 = v$RD_5912_out0 && v$RM_11352_out0;
assign v$G2_12767_out0 = v$RD_6376_out0 && v$RM_11816_out0;
assign v$TX$inst0_608_out0 = v$TX$INSTUCTION0_228_out0;
assign v$MUX1_1735_out0 = v$EXEC1_20_out0 ? v$RMN_13437_out0 : v$RAMDOUT_2414_out0;
assign v$MUX1_1736_out0 = v$EXEC1_21_out0 ? v$RMN_13438_out0 : v$RAMDOUT_2415_out0;
assign v$CARRY_4912_out0 = v$G2_12303_out0;
assign v$CARRY_5376_out0 = v$G2_12767_out0;
assign v$RX$INSTRUCTION_8686_out0 = v$RX$INST_2334_out0;
assign v$RD$SIG$NEW_8759_out0 = v$MUX2_188_out0;
assign v$RD$SIG$NEW_8760_out0 = v$MUX2_189_out0;
assign v$S_8913_out0 = v$G1_7767_out0;
assign v$S_9377_out0 = v$G1_8231_out0;
assign v$_10536_out0 = v$IN_2350_out0[15:15];
assign v$_10537_out0 = v$IN_2351_out0[15:15];
assign v$OP2$SIG$NEW_11190_out0 = v$MUX1_7702_out0;
assign v$OP2$SIG$NEW_11191_out0 = v$MUX1_7703_out0;
assign v$_13291_out0 = v$IN_2350_out0[3:0];
assign v$_13291_out1 = v$IN_2350_out0[15:12];
assign v$_13292_out0 = v$IN_2351_out0[3:0];
assign v$_13292_out1 = v$IN_2351_out0[15:12];
assign v$_164_out0 = { v$_13291_out1,v$_10536_out0 };
assign v$_165_out0 = { v$_13292_out1,v$_10537_out0 };
assign v$S_1242_out0 = v$S_8913_out0;
assign v$S_1466_out0 = v$S_9377_out0;
assign v$G1_4018_out0 = v$CARRY_4912_out0 || v$CARRY_4911_out0;
assign v$G1_4242_out0 = v$CARRY_5376_out0 || v$CARRY_5375_out0;
assign v$RX$INSTRUCTION_4659_out0 = v$RX$INSTRUCTION_8686_out0;
assign v$MUX5_7678_out0 = v$TX$inst0_608_out0 ? v$BYTE$COMP$10_13611_out0 : v$BYTE$COMP$11_1163_out0;
assign v$RD$SIG$NEW_10872_out0 = v$RD$SIG$NEW_8759_out0;
assign v$RD$SIG$NEW_10873_out0 = v$RD$SIG$NEW_8760_out0;
assign v$REGDIN_11041_out0 = v$MUX1_1735_out0;
assign v$REGDIN_11042_out0 = v$MUX1_1736_out0;
assign v$OP2$SIG$NEW_11218_out0 = v$OP2$SIG$NEW_11190_out0;
assign v$OP2$SIG$NEW_11219_out0 = v$OP2$SIG$NEW_11191_out0;
assign v$NOTUSED_13265_out0 = v$_13291_out0;
assign v$NOTUSED_13266_out0 = v$_13292_out0;
assign v$G22_13663_out0 = v$TX$inst0_608_out0 || v$TX$INSTUCTION1_4859_out0;
assign v$RD$SIG_109_out0 = v$RD$SIG$NEW_10872_out0;
assign v$RD$SIG_110_out0 = v$RD$SIG$NEW_10873_out0;
assign v$COUT_710_out0 = v$G1_4018_out0;
assign v$COUT_934_out0 = v$G1_4242_out0;
assign v$_2553_out0 = { v$_4783_out0,v$S_1242_out0 };
assign v$_2568_out0 = { v$_4798_out0,v$S_1466_out0 };
assign v$LS$REGIN_3303_out0 = v$REGDIN_11041_out0;
assign v$LS$REGIN_3304_out0 = v$REGDIN_11042_out0;
assign v$byte$comp$1_6923_out0 = v$MUX5_7678_out0;
assign v$_11055_out0 = { v$_164_out0,v$_10536_out0 };
assign v$_11056_out0 = { v$_165_out0,v$_10537_out0 };
assign v$TX$INST_11239_out0 = v$G22_13663_out0;
assign v$OP2$SIG_13314_out0 = v$OP2$SIG$NEW_11218_out0;
assign v$OP2$SIG_13315_out0 = v$OP2$SIG$NEW_11219_out0;
assign v$RX$INSTRUCTION_13325_out0 = v$RX$INSTRUCTION_4659_out0;
assign v$_3178_out0 = { v$OP2$SIG_13314_out0,v$C4_2593_out0 };
assign v$_3179_out0 = { v$OP2$SIG_13315_out0,v$C4_2594_out0 };
assign v$byte$comp$1_6872_out0 = v$byte$comp$1_6923_out0;
assign v$G4_6915_out0 = ! v$RX$INSTRUCTION_13325_out0;
assign v$G8_7103_out0 = v$RX$INSTRUCTION_13325_out0 || v$RXBYTERECEIVED_3269_out0;
assign v$CIN_9826_out0 = v$COUT_710_out0;
assign v$CIN_10050_out0 = v$COUT_934_out0;
assign v$G18_10489_out0 = ! v$RX$INSTRUCTION_13325_out0;
assign v$TX$INSTRUCTION_10501_out0 = v$TX$INST_11239_out0;
assign v$_11231_out0 = { v$_11055_out0,v$_10536_out0 };
assign v$_11232_out0 = { v$_11056_out0,v$_10537_out0 };
assign v$_13275_out0 = { v$RD$SIG_109_out0,v$C4_2593_out0 };
assign v$_13276_out0 = { v$RD$SIG_110_out0,v$C4_2594_out0 };
assign v$_2791_out0 = { v$_11231_out0,v$_10536_out0 };
assign v$_2792_out0 = { v$_11232_out0,v$_10537_out0 };
assign v$G3_3948_out0 = v$G4_6915_out0 && v$G1_10476_out0;
assign v$XOR2_4486_out0 = v$_3178_out0 ^ v$C11_4539_out0;
assign v$XOR2_4487_out0 = v$_3179_out0 ^ v$C11_4540_out0;
assign v$RD_5900_out0 = v$CIN_9826_out0;
assign v$RD_6364_out0 = v$CIN_10050_out0;
assign v$G16_7701_out0 = v$G19_3860_out0 && v$G18_10489_out0;
assign v$BYTE$COMP$1_8743_out0 = v$byte$comp$1_6872_out0;
assign v$XOR1_11246_out0 = v$_13275_out0 ^ v$C5_2688_out0;
assign v$XOR1_11247_out0 = v$_13276_out0 ^ v$C5_2689_out0;
assign v$TX$INSTRUCTION_13631_out0 = v$TX$INSTRUCTION_10501_out0;
assign v$OUT_460_out0 = v$_2791_out0;
assign v$OUT_461_out0 = v$_2792_out0;
assign {v$A5_1901_out1,v$A5_1901_out0 } = v$C7_1865_out0 + v$XOR2_4486_out0 + v$C12_1151_out0;
assign {v$A5_1902_out1,v$A5_1902_out0 } = v$C7_1866_out0 + v$XOR2_4487_out0 + v$C12_1152_out0;
assign v$TX$INSTRUCTION_6875_out0 = v$TX$INSTRUCTION_13631_out0;
assign v$G1_7755_out0 = ((v$RD_5900_out0 && !v$RM_11340_out0) || (!v$RD_5900_out0) && v$RM_11340_out0);
assign v$G1_8219_out0 = ((v$RD_6364_out0 && !v$RM_11804_out0) || (!v$RD_6364_out0) && v$RM_11804_out0);
assign v$G5_10801_out0 = v$G3_3948_out0 && v$_2983_out0;
assign v$G20_11040_out0 = v$G17_1903_out0 || v$G16_7701_out0;
assign v$G7_11095_out0 = v$G6_4818_out0 && v$G3_3948_out0;
assign {v$A4_11227_out1,v$A4_11227_out0 } = v$XOR1_11246_out0 + v$C7_1865_out0 + v$C6_10317_out0;
assign {v$A4_11228_out1,v$A4_11228_out0 } = v$XOR1_11247_out0 + v$C7_1866_out0 + v$C6_10318_out0;
assign v$G2_12291_out0 = v$RD_5900_out0 && v$RM_11340_out0;
assign v$G2_12755_out0 = v$RD_6364_out0 && v$RM_11804_out0;
assign v$TX$INSTRUCTION_453_out0 = v$TX$INSTRUCTION_6875_out0;
assign v$MUX2_1181_out0 = v$G1_289_out0 ? v$A5_1901_out0 : v$_3178_out0;
assign v$MUX2_1182_out0 = v$G1_290_out0 ? v$A5_1902_out0 : v$_3179_out0;
assign v$MUX1_1883_out0 = v$RD$SIGN_2405_out0 ? v$A4_11227_out0 : v$_13275_out0;
assign v$MUX1_1884_out0 = v$RD$SIGN_2406_out0 ? v$A4_11228_out0 : v$_13276_out0;
assign v$MUX3_3041_out0 = v$ASR_10566_out0 ? v$OUT_460_out0 : v$MUX2_13319_out0;
assign v$MUX3_3042_out0 = v$ASR_10567_out0 ? v$OUT_461_out0 : v$MUX2_13320_out0;
assign v$CARRY_4900_out0 = v$G2_12291_out0;
assign v$CARRY_5364_out0 = v$G2_12755_out0;
assign v$S_8901_out0 = v$G1_7755_out0;
assign v$S_9365_out0 = v$G1_8219_out0;
assign v$NOTUSED4_10530_out0 = v$A4_11227_out1;
assign v$NOTUSED4_10531_out0 = v$A4_11228_out1;
assign v$NOTUSED1_10684_out0 = v$A5_1901_out1;
assign v$NOTUSED1_10685_out0 = v$A5_1902_out1;
assign v$G10_10694_out0 = v$G5_10801_out0 || v$G9_13655_out0;
assign v$S_1237_out0 = v$S_8901_out0;
assign v$S_1461_out0 = v$S_9365_out0;
assign v$TRANSMIT$INSTRUCTION_1713_out0 = v$TX$INSTRUCTION_453_out0;
assign v$TX$INSTRUCTION_2825_out0 = v$TX$INSTRUCTION_453_out0;
assign v$G1_4013_out0 = v$CARRY_4900_out0 || v$CARRY_4899_out0;
assign v$G1_4237_out0 = v$CARRY_5364_out0 || v$CARRY_5363_out0;
assign v$_4488_out0 = v$MUX3_3041_out0[3:0];
assign v$_4488_out1 = v$MUX3_3041_out0[15:12];
assign v$_4489_out0 = v$MUX3_3042_out0[3:0];
assign v$_4489_out1 = v$MUX3_3042_out0[15:12];
assign v$_4547_out0 = { v$G7_11095_out0,v$G10_10694_out0 };
assign {v$A6_10463_out1,v$A6_10463_out0 } = v$MUX1_1883_out0 + v$MUX2_1181_out0 + v$C3_4741_out0;
assign {v$A6_10464_out1,v$A6_10464_out0 } = v$MUX1_1884_out0 + v$MUX2_1182_out0 + v$C3_4742_out0;
assign v$_167_out0 = { v$_4488_out1,v$_4488_out0 };
assign v$_168_out0 = { v$_4489_out1,v$_4489_out0 };
assign v$COUT_705_out0 = v$G1_4013_out0;
assign v$COUT_929_out0 = v$G1_4237_out0;
assign v$SEL1_2305_out0 = v$A6_10463_out0[15:15];
assign v$SEL1_2306_out0 = v$A6_10464_out0[15:15];
assign v$G23_2614_out0 = v$G21_10681_out0 && v$TX$INSTRUCTION_2825_out0;
assign v$transmit$INSTRUCTION_2674_out0 = v$TRANSMIT$INSTRUCTION_1713_out0;
assign v$_7033_out0 = { v$_2553_out0,v$S_1237_out0 };
assign v$_7048_out0 = { v$_2568_out0,v$S_1461_out0 };
assign v$NOTUSED_10835_out0 = v$A6_10463_out1;
assign v$NOTUSED_10836_out0 = v$A6_10464_out1;
assign v$MUX1_11061_out0 = v$RX$INSTRUCTION_13325_out0 ? v$C5_10356_out0 : v$_4547_out0;
assign v$XOR3_13599_out0 = v$A6_10463_out0 ^ v$C15_1730_out0;
assign v$XOR3_13600_out0 = v$A6_10464_out0 ^ v$C15_1731_out0;
assign v$SIGN$ANS_1970_out0 = v$SEL1_2305_out0;
assign v$SIGN$ANS_1971_out0 = v$SEL1_2306_out0;
assign v$MUX4_2229_out0 = v$ROR_544_out0 ? v$_167_out0 : v$MUX3_3041_out0;
assign v$MUX4_2230_out0 = v$ROR_545_out0 ? v$_168_out0 : v$MUX3_3042_out0;
assign v$MUX8_2697_out0 = v$transmit$INSTRUCTION_2674_out0 ? v$C1_10259_out0 : v$FF8_11222_out0;
assign v$CIN_9825_out0 = v$COUT_705_out0;
assign v$CIN_10049_out0 = v$COUT_929_out0;
assign v$G24_10460_out0 = ! v$G23_2614_out0;
assign v$G2_10471_out0 = ! v$transmit$INSTRUCTION_2674_out0;
assign v$MUX3_10994_out0 = v$G25_4658_out0 ? v$G23_2614_out0 : v$C7_3222_out0;
assign {v$A8_11155_out1,v$A8_11155_out0 } = v$XOR3_13599_out0 + v$C13_2185_out0 + v$C14_1674_out0;
assign {v$A8_11156_out1,v$A8_11156_out0 } = v$XOR3_13600_out0 + v$C13_2186_out0 + v$C14_1675_out0;
assign v$G3_13507_out0 = v$transmit$INSTRUCTION_2674_out0 || v$SHIFHT$ENABLE_13501_out0;
assign v$TX$OVERFLOW_500_out0 = v$MUX3_10994_out0;
assign v$G10_602_out0 = v$G7_2455_out0 && v$G2_10471_out0;
assign v$_1813_out0 = { v$MUX3_10994_out0,v$C4_1201_out0 };
assign v$ENABLE_2651_out0 = v$G3_13507_out0;
assign v$NOTUSED2_5794_out0 = v$A8_11155_out1;
assign v$NOTUSED2_5795_out0 = v$A8_11156_out1;
assign v$RD_5898_out0 = v$CIN_9825_out0;
assign v$RD_6362_out0 = v$CIN_10049_out0;
assign v$STARTBIT_6968_out0 = v$G2_10471_out0;
assign v$STARTBIT_6970_out0 = v$G24_10460_out0;
assign v$SIGN$ANS_8650_out0 = v$SIGN$ANS_1970_out0;
assign v$SIGN$ANS_8651_out0 = v$SIGN$ANS_1971_out0;
assign v$MUX3_8669_out0 = v$SEL1_2305_out0 ? v$A8_11155_out0 : v$A6_10463_out0;
assign v$MUX3_8670_out0 = v$SEL1_2306_out0 ? v$A8_11156_out0 : v$A6_10464_out0;
assign v$MUX5_10605_out0 = v$EN_13181_out0 ? v$MUX4_2229_out0 : v$IN_13548_out0;
assign v$MUX5_10606_out0 = v$EN_13182_out0 ? v$MUX4_2230_out0 : v$IN_13549_out0;
assign v$MUX9_166_out0 = v$G10_602_out0 ? v$2_7072_out0 : v$FF9_8805_out0;
assign v$OUT_2352_out0 = v$MUX5_10605_out0;
assign v$OUT_2353_out0 = v$MUX5_10606_out0;
assign v$SIGN$ANS_4457_out0 = v$SIGN$ANS_8650_out0;
assign v$SIGN$ANS_4458_out0 = v$SIGN$ANS_8651_out0;
assign v$G1_7753_out0 = ((v$RD_5898_out0 && !v$RM_11338_out0) || (!v$RD_5898_out0) && v$RM_11338_out0);
assign v$G1_8217_out0 = ((v$RD_6362_out0 && !v$RM_11802_out0) || (!v$RD_6362_out0) && v$RM_11802_out0);
assign v$G35_10361_out0 = v$STARTBIT_6968_out0 && v$G36_3136_out0;
assign v$G35_10363_out0 = v$STARTBIT_6970_out0 && v$G36_3138_out0;
assign v$TX$OVERFLOW_10481_out0 = v$TX$OVERFLOW_500_out0;
assign v$SEL8_10686_out0 = v$MUX3_8669_out0[11:0];
assign v$SEL8_10687_out0 = v$MUX3_8670_out0[11:0];
assign v$G2_12289_out0 = v$RD_5898_out0 && v$RM_11338_out0;
assign v$G2_12753_out0 = v$RD_6362_out0 && v$RM_11802_out0;
assign v$IN_190_out0 = v$OUT_2352_out0;
assign v$IN_191_out0 = v$OUT_2353_out0;
assign v$ENABLE_2019_out0 = v$G35_10361_out0;
assign v$ENABLE_2021_out0 = v$G35_10363_out0;
assign v$OUTSTREAM_2097_out0 = v$MUX9_166_out0;
assign v$CARRY_4898_out0 = v$G2_12289_out0;
assign v$CARRY_5362_out0 = v$G2_12753_out0;
assign v$S_8899_out0 = v$G1_7753_out0;
assign v$S_9363_out0 = v$G1_8217_out0;
assign v$SIGN$ANS_10302_out0 = v$SIGN$ANS_4457_out0;
assign v$SIGN$ANS_10303_out0 = v$SIGN$ANS_4458_out0;
assign v$TX$OVERFLOW_13294_out0 = v$TX$OVERFLOW_10481_out0;
assign v$OUT_22_out0 = v$OUTSTREAM_2097_out0;
assign v$IN_685_out0 = v$IN_190_out0;
assign v$IN_686_out0 = v$IN_191_out0;
assign v$S_1236_out0 = v$S_8899_out0;
assign v$S_1460_out0 = v$S_9363_out0;
assign v$_3125_out0 = v$IN_190_out0[7:0];
assign v$_3125_out1 = v$IN_190_out0[15:8];
assign v$_3126_out0 = v$IN_191_out0[7:0];
assign v$_3126_out1 = v$IN_191_out0[15:8];
assign v$G1_4012_out0 = v$CARRY_4898_out0 || v$CARRY_4897_out0;
assign v$G1_4236_out0 = v$CARRY_5362_out0 || v$CARRY_5361_out0;
assign v$G18_8800_out0 = !(v$ENABLE_2019_out0 || v$Q7_6889_out0);
assign v$G18_8802_out0 = !(v$ENABLE_2021_out0 || v$Q7_6891_out0);
assign v$NOTUSED2_41_out0 = v$_3125_out1;
assign v$NOTUSED2_42_out0 = v$_3126_out1;
assign v$COUT_704_out0 = v$G1_4012_out0;
assign v$COUT_928_out0 = v$G1_4236_out0;
assign v$BIT$OUT_2015_out0 = v$OUT_22_out0;
assign v$G21_3809_out0 = v$G18_8800_out0 || v$G22_10984_out0;
assign v$G21_3811_out0 = v$G18_8802_out0 || v$G22_10986_out0;
assign v$_4709_out0 = { v$C1_13446_out0,v$_3125_out0 };
assign v$_4710_out0 = { v$C1_13447_out0,v$_3126_out0 };
assign v$_13519_out0 = { v$_7033_out0,v$S_1236_out0 };
assign v$_13534_out0 = { v$_7048_out0,v$S_1460_out0 };
assign v$BIT_383_out0 = v$BIT$OUT_2015_out0;
assign v$CIN_9832_out0 = v$COUT_704_out0;
assign v$CIN_10056_out0 = v$COUT_928_out0;
assign v$MUX1_10443_out0 = v$LSL_1861_out0 ? v$_4709_out0 : v$IN_685_out0;
assign v$MUX1_10444_out0 = v$LSL_1862_out0 ? v$_4710_out0 : v$IN_686_out0;
assign v$BIT$OUT_10705_out0 = v$BIT$OUT_2015_out0;
assign v$G2_3214_out0 = ! v$BIT_383_out0;
assign v$RD_5914_out0 = v$CIN_9832_out0;
assign v$RD_6378_out0 = v$CIN_10056_out0;
assign v$STARTBIT_6969_out0 = v$BIT_383_out0;
assign v$_8673_out0 = v$MUX1_10443_out0[7:0];
assign v$_8673_out1 = v$MUX1_10443_out0[15:8];
assign v$_8674_out0 = v$MUX1_10444_out0[7:0];
assign v$_8674_out1 = v$MUX1_10444_out0[15:8];
assign v$BIT$OUT_13326_out0 = v$BIT$OUT_10705_out0;
assign v$MUX2_1180_out0 = v$G22_10620_out0 ? v$G2_3214_out0 : v$C6_1732_out0;
assign v$G1_7769_out0 = ((v$RD_5914_out0 && !v$RM_11354_out0) || (!v$RD_5914_out0) && v$RM_11354_out0);
assign v$G1_8233_out0 = ((v$RD_6378_out0 && !v$RM_11818_out0) || (!v$RD_6378_out0) && v$RM_11818_out0);
assign v$G35_10362_out0 = v$STARTBIT_6969_out0 && v$G36_3137_out0;
assign v$_10504_out0 = { v$_8673_out1,v$C1_13446_out0 };
assign v$_10505_out0 = { v$_8674_out1,v$C1_13447_out0 };
assign v$NOTUSED_10564_out0 = v$_8673_out0;
assign v$NOTUSED_10565_out0 = v$_8674_out0;
assign v$G2_12305_out0 = v$RD_5914_out0 && v$RM_11354_out0;
assign v$G2_12769_out0 = v$RD_6378_out0 && v$RM_11818_out0;
assign v$ENABLE_2020_out0 = v$G35_10362_out0;
assign v$MUX2_2337_out0 = v$LSR_1174_out0 ? v$_10504_out0 : v$MUX1_10443_out0;
assign v$MUX2_2338_out0 = v$LSR_1175_out0 ? v$_10505_out0 : v$MUX1_10444_out0;
assign v$CARRY_4914_out0 = v$G2_12305_out0;
assign v$CARRY_5378_out0 = v$G2_12769_out0;
assign v$TX$PROGRESS_8645_out0 = v$MUX2_1180_out0;
assign v$S_8915_out0 = v$G1_7769_out0;
assign v$S_9379_out0 = v$G1_8233_out0;
assign v$_13337_out0 = { v$MUX2_1180_out0,v$C3_10853_out0 };
assign v$TX$IN$PROGRESS_235_out0 = v$TX$PROGRESS_8645_out0;
assign v$S_1243_out0 = v$S_8915_out0;
assign v$S_1467_out0 = v$S_9379_out0;
assign v$_2425_out0 = { v$_13337_out0,v$_1813_out0 };
assign v$G1_4019_out0 = v$CARRY_4914_out0 || v$CARRY_4913_out0;
assign v$G1_4243_out0 = v$CARRY_5378_out0 || v$CARRY_5377_out0;
assign v$IN_5796_out0 = v$MUX2_2337_out0;
assign v$IN_5797_out0 = v$MUX2_2338_out0;
assign v$G18_8801_out0 = !(v$ENABLE_2020_out0 || v$Q7_6890_out0);
assign v$COUT_711_out0 = v$G1_4019_out0;
assign v$COUT_935_out0 = v$G1_4243_out0;
assign v$_2582_out0 = v$IN_5796_out0[7:0];
assign v$_2582_out1 = v$IN_5796_out0[15:8];
assign v$_2583_out0 = v$IN_5797_out0[7:0];
assign v$_2583_out1 = v$IN_5797_out0[15:8];
assign v$_3266_out0 = v$IN_5796_out0[15:15];
assign v$_3267_out0 = v$IN_5797_out0[15:15];
assign v$_3312_out0 = { v$_13519_out0,v$S_1243_out0 };
assign v$_3327_out0 = { v$_13534_out0,v$S_1467_out0 };
assign v$G21_3810_out0 = v$G18_8801_out0 || v$G22_10985_out0;
assign v$_10532_out0 = { v$_10376_out0,v$_2425_out0 };
assign v$TX$IN$PROGRESS_13634_out0 = v$TX$IN$PROGRESS_235_out0;
assign v$NOTUSED_68_out0 = v$_2582_out0;
assign v$NOTUSED_69_out0 = v$_2583_out0;
assign v$_7704_out0 = { v$_2582_out1,v$_3266_out0 };
assign v$_7705_out0 = { v$_2583_out1,v$_3267_out0 };
assign v$CIN_9833_out0 = v$COUT_711_out0;
assign v$CIN_10057_out0 = v$COUT_935_out0;
assign v$RD$STATUS_10500_out0 = v$_10532_out0;
assign v$RD_5916_out0 = v$CIN_9833_out0;
assign v$RD_6380_out0 = v$CIN_10057_out0;
assign v$STATUS$REGISTER_10359_out0 = v$RD$STATUS_10500_out0;
assign v$_10806_out0 = { v$_7704_out0,v$_3266_out0 };
assign v$_10807_out0 = { v$_7705_out0,v$_3267_out0 };
assign v$STATUS$REGISTER_185_out0 = v$STATUS$REGISTER_10359_out0;
assign v$G1_7771_out0 = ((v$RD_5916_out0 && !v$RM_11356_out0) || (!v$RD_5916_out0) && v$RM_11356_out0);
assign v$G1_8235_out0 = ((v$RD_6380_out0 && !v$RM_11820_out0) || (!v$RD_6380_out0) && v$RM_11820_out0);
assign v$G2_12307_out0 = v$RD_5916_out0 && v$RM_11356_out0;
assign v$G2_12771_out0 = v$RD_6380_out0 && v$RM_11820_out0;
assign v$_13310_out0 = { v$_10806_out0,v$_3266_out0 };
assign v$_13311_out0 = { v$_10807_out0,v$_3267_out0 };
assign v$_107_out0 = { v$_13310_out0,v$_3266_out0 };
assign v$_108_out0 = { v$_13311_out0,v$_3267_out0 };
assign v$CARRY_4916_out0 = v$G2_12307_out0;
assign v$CARRY_5380_out0 = v$G2_12771_out0;
assign v$S_8917_out0 = v$G1_7771_out0;
assign v$S_9381_out0 = v$G1_8235_out0;
assign v$STATUS$REGISTER_13778_out0 = v$STATUS$REGISTER_185_out0;
assign v$S_1244_out0 = v$S_8917_out0;
assign v$S_1468_out0 = v$S_9381_out0;
assign v$STATUS$REGISTER_2866_out0 = v$STATUS$REGISTER_13778_out0;
assign v$STATUS$REGISTER_2867_out0 = v$STATUS$REGISTER_13778_out0;
assign v$G1_4020_out0 = v$CARRY_4916_out0 || v$CARRY_4915_out0;
assign v$G1_4244_out0 = v$CARRY_5380_out0 || v$CARRY_5379_out0;
assign v$_5851_out0 = { v$_107_out0,v$_3266_out0 };
assign v$_5852_out0 = { v$_108_out0,v$_3267_out0 };
assign v$_538_out0 = { v$_5851_out0,v$_3266_out0 };
assign v$_539_out0 = { v$_5852_out0,v$_3267_out0 };
assign v$COUT_712_out0 = v$G1_4020_out0;
assign v$COUT_936_out0 = v$G1_4244_out0;
assign v$STATUS$REGISTER_5858_out0 = v$STATUS$REGISTER_2866_out0;
assign v$STATUS$REGISTER_5859_out0 = v$STATUS$REGISTER_2867_out0;
assign v$_7148_out0 = { v$_3312_out0,v$S_1244_out0 };
assign v$_7163_out0 = { v$_3327_out0,v$S_1468_out0 };
assign v$_2223_out0 = { v$_538_out0,v$_3266_out0 };
assign v$_2224_out0 = { v$_539_out0,v$_3267_out0 };
assign v$MUX4_4579_out0 = v$STAT$INSTRUCTION_2855_out0 ? v$STATUS$REGISTER_5858_out0 : v$RAM$OUT_11214_out0;
assign v$MUX4_4580_out0 = v$STAT$INSTRUCTION_2856_out0 ? v$STATUS$REGISTER_5859_out0 : v$RAM$OUT_11215_out0;
assign v$CIN_9835_out0 = v$COUT_712_out0;
assign v$CIN_10059_out0 = v$COUT_936_out0;
assign v$DFQDF_3025_out0 = v$MUX4_4579_out0;
assign v$DFQDF_3026_out0 = v$MUX4_4580_out0;
assign v$RD_5920_out0 = v$CIN_9835_out0;
assign v$RD_6384_out0 = v$CIN_10059_out0;
assign v$_7124_out0 = { v$_2223_out0,v$_3266_out0 };
assign v$_7125_out0 = { v$_2224_out0,v$_3267_out0 };
assign v$OUT_2857_out0 = v$_7124_out0;
assign v$OUT_2858_out0 = v$_7125_out0;
assign v$G1_7775_out0 = ((v$RD_5920_out0 && !v$RM_11360_out0) || (!v$RD_5920_out0) && v$RM_11360_out0);
assign v$G1_8239_out0 = ((v$RD_6384_out0 && !v$RM_11824_out0) || (!v$RD_6384_out0) && v$RM_11824_out0);
assign v$G2_12311_out0 = v$RD_5920_out0 && v$RM_11360_out0;
assign v$G2_12775_out0 = v$RD_6384_out0 && v$RM_11824_out0;
assign v$CARRY_4920_out0 = v$G2_12311_out0;
assign v$CARRY_5384_out0 = v$G2_12775_out0;
assign v$MUX3_6864_out0 = v$ASR_10366_out0 ? v$OUT_2857_out0 : v$MUX2_2337_out0;
assign v$MUX3_6865_out0 = v$ASR_10367_out0 ? v$OUT_2858_out0 : v$MUX2_2338_out0;
assign v$S_8921_out0 = v$G1_7775_out0;
assign v$S_9385_out0 = v$G1_8239_out0;
assign v$S_1246_out0 = v$S_8921_out0;
assign v$S_1470_out0 = v$S_9385_out0;
assign v$G1_4022_out0 = v$CARRY_4920_out0 || v$CARRY_4919_out0;
assign v$G1_4246_out0 = v$CARRY_5384_out0 || v$CARRY_5383_out0;
assign v$_11132_out0 = v$MUX3_6864_out0[7:0];
assign v$_11132_out1 = v$MUX3_6864_out0[15:8];
assign v$_11133_out0 = v$MUX3_6865_out0[7:0];
assign v$_11133_out1 = v$MUX3_6865_out0[15:8];
assign v$COUT_714_out0 = v$G1_4022_out0;
assign v$COUT_938_out0 = v$G1_4246_out0;
assign v$_4750_out0 = { v$_7148_out0,v$S_1246_out0 };
assign v$_4765_out0 = { v$_7163_out0,v$S_1470_out0 };
assign v$_6870_out0 = { v$_11132_out1,v$_11132_out0 };
assign v$_6871_out0 = { v$_11133_out1,v$_11133_out0 };
assign v$CIN_9828_out0 = v$COUT_714_out0;
assign v$CIN_10052_out0 = v$COUT_938_out0;
assign v$MUX4_13498_out0 = v$ROR_282_out0 ? v$_6870_out0 : v$MUX3_6864_out0;
assign v$MUX4_13499_out0 = v$ROR_283_out0 ? v$_6871_out0 : v$MUX3_6865_out0;
assign v$MUX5_3305_out0 = v$EN_2445_out0 ? v$MUX4_13498_out0 : v$IN_685_out0;
assign v$MUX5_3306_out0 = v$EN_2446_out0 ? v$MUX4_13499_out0 : v$IN_686_out0;
assign v$RD_5906_out0 = v$CIN_9828_out0;
assign v$RD_6370_out0 = v$CIN_10052_out0;
assign v$G1_7761_out0 = ((v$RD_5906_out0 && !v$RM_11346_out0) || (!v$RD_5906_out0) && v$RM_11346_out0);
assign v$G1_8225_out0 = ((v$RD_6370_out0 && !v$RM_11810_out0) || (!v$RD_6370_out0) && v$RM_11810_out0);
assign v$OUT_10264_out0 = v$MUX5_3305_out0;
assign v$OUT_10265_out0 = v$MUX5_3306_out0;
assign v$G2_12297_out0 = v$RD_5906_out0 && v$RM_11346_out0;
assign v$G2_12761_out0 = v$RD_6370_out0 && v$RM_11810_out0;
assign v$OP2_2862_out0 = v$OUT_10264_out0;
assign v$OP2_2863_out0 = v$OUT_10265_out0;
assign v$CARRY_4906_out0 = v$G2_12297_out0;
assign v$CARRY_5370_out0 = v$G2_12761_out0;
assign v$S_8907_out0 = v$G1_7761_out0;
assign v$S_9371_out0 = v$G1_8225_out0;
assign v$S_1239_out0 = v$S_8907_out0;
assign v$S_1463_out0 = v$S_9371_out0;
assign v$G1_4015_out0 = v$CARRY_4906_out0 || v$CARRY_4905_out0;
assign v$G1_4239_out0 = v$CARRY_5370_out0 || v$CARRY_5369_out0;
assign v$OP2_11153_out0 = v$OP2_2862_out0;
assign v$OP2_11154_out0 = v$OP2_2863_out0;
assign v$COUT_707_out0 = v$G1_4015_out0;
assign v$COUT_931_out0 = v$G1_4239_out0;
assign v$OP2_3940_out0 = v$OP2_11153_out0;
assign v$OP2_3941_out0 = v$OP2_11154_out0;
assign v$_6927_out0 = { v$_4750_out0,v$S_1239_out0 };
assign v$_6942_out0 = { v$_4765_out0,v$S_1463_out0 };
assign v$OP2_2322_out0 = v$OP2_3940_out0;
assign v$OP2_2323_out0 = v$OP2_3941_out0;
assign v$CIN_9829_out0 = v$COUT_707_out0;
assign v$CIN_10053_out0 = v$COUT_931_out0;
assign v$RD_5908_out0 = v$CIN_9829_out0;
assign v$RD_6372_out0 = v$CIN_10053_out0;
assign v$OP2_10751_out0 = v$OP2_2322_out0;
assign v$OP2_10752_out0 = v$OP2_2323_out0;
assign v$MUX5_2595_out0 = v$MOV_196_out0 ? v$OP2_10751_out0 : v$OP1_2060_out0;
assign v$MUX5_2596_out0 = v$MOV_197_out0 ? v$OP2_10752_out0 : v$OP1_2061_out0;
assign v$B_3350_out0 = v$OP2_10751_out0;
assign v$B_3352_out0 = v$OP2_10752_out0;
assign v$G1_7763_out0 = ((v$RD_5908_out0 && !v$RM_11348_out0) || (!v$RD_5908_out0) && v$RM_11348_out0);
assign v$G1_8227_out0 = ((v$RD_6372_out0 && !v$RM_11812_out0) || (!v$RD_6372_out0) && v$RM_11812_out0);
assign v$A_11250_out0 = v$OP2_10751_out0;
assign v$A_11252_out0 = v$OP2_10752_out0;
assign v$G2_12299_out0 = v$RD_5908_out0 && v$RM_11348_out0;
assign v$G2_12763_out0 = v$RD_6372_out0 && v$RM_11812_out0;
assign v$_77_out0 = v$A_11250_out0[3:3];
assign v$_79_out0 = v$A_11252_out0[3:3];
assign v$_192_out0 = v$A_11250_out0[15:15];
assign v$_194_out0 = v$A_11252_out0[15:15];
assign v$_198_out0 = v$B_3350_out0[7:7];
assign v$_199_out0 = v$B_3352_out0[7:7];
assign v$_321_out0 = v$A_11250_out0[0:0];
assign v$_323_out0 = v$A_11252_out0[0:0];
assign v$_329_out0 = v$A_11250_out0[9:9];
assign v$_331_out0 = v$A_11252_out0[9:9];
assign v$_1722_out0 = v$B_3350_out0[5:5];
assign v$_1723_out0 = v$B_3352_out0[5:5];
assign v$_1904_out0 = v$B_3350_out0[9:9];
assign v$_1905_out0 = v$B_3352_out0[9:9];
assign v$_2093_out0 = v$A_11250_out0[13:13];
assign v$_2095_out0 = v$A_11252_out0[13:13];
assign v$_2418_out0 = v$A_11250_out0[6:6];
assign v$_2420_out0 = v$A_11252_out0[6:6];
assign v$_2462_out0 = v$B_3350_out0[2:2];
assign v$_2463_out0 = v$B_3352_out0[2:2];
assign v$_2943_out0 = v$B_3350_out0[10:10];
assign v$_2944_out0 = v$B_3352_out0[10:10];
assign v$_3119_out0 = v$A_11250_out0[14:14];
assign v$_3121_out0 = v$A_11252_out0[14:14];
assign v$_3237_out0 = v$B_3350_out0[11:11];
assign v$_3238_out0 = v$B_3352_out0[11:11];
assign v$_3282_out0 = v$A_11250_out0[2:2];
assign v$_3284_out0 = v$A_11252_out0[2:2];
assign v$_4610_out0 = v$B_3350_out0[3:3];
assign v$_4611_out0 = v$B_3352_out0[3:3];
assign v$_4812_out0 = v$B_3350_out0[4:4];
assign v$_4813_out0 = v$B_3352_out0[4:4];
assign v$_4814_out0 = v$B_3350_out0[14:14];
assign v$_4815_out0 = v$B_3352_out0[14:14];
assign v$_4833_out0 = v$B_3350_out0[6:6];
assign v$_4834_out0 = v$B_3352_out0[6:6];
assign v$CARRY_4908_out0 = v$G2_12299_out0;
assign v$CARRY_5372_out0 = v$G2_12763_out0;
assign v$_7070_out0 = v$B_3350_out0[0:0];
assign v$_7071_out0 = v$B_3352_out0[0:0];
assign v$_8748_out0 = v$A_11250_out0[8:8];
assign v$_8750_out0 = v$A_11252_out0[8:8];
assign v$_8827_out0 = v$A_11250_out0[7:7];
assign v$_8829_out0 = v$A_11252_out0[7:7];
assign v$_8831_out0 = v$B_3350_out0[15:15];
assign v$_8832_out0 = v$B_3352_out0[15:15];
assign v$S_8909_out0 = v$G1_7763_out0;
assign v$S_9373_out0 = v$G1_8227_out0;
assign v$_10377_out0 = v$A_11250_out0[5:5];
assign v$_10379_out0 = v$A_11252_out0[5:5];
assign v$_10385_out0 = v$A_11250_out0[1:1];
assign v$_10387_out0 = v$A_11252_out0[1:1];
assign v$_10538_out0 = v$B_3350_out0[13:13];
assign v$_10539_out0 = v$B_3352_out0[13:13];
assign v$_10695_out0 = v$A_11250_out0[4:4];
assign v$_10697_out0 = v$A_11252_out0[4:4];
assign v$_10777_out0 = v$A_11250_out0[12:12];
assign v$_10779_out0 = v$A_11252_out0[12:12];
assign v$_10862_out0 = v$A_11250_out0[10:10];
assign v$_10864_out0 = v$A_11252_out0[10:10];
assign v$_11212_out0 = v$B_3350_out0[12:12];
assign v$_11213_out0 = v$B_3352_out0[12:12];
assign v$_13251_out0 = v$B_3350_out0[1:1];
assign v$_13252_out0 = v$B_3352_out0[1:1];
assign v$_13392_out0 = v$B_3350_out0[8:8];
assign v$_13393_out0 = v$B_3352_out0[8:8];
assign v$_13552_out0 = v$A_11250_out0[11:11];
assign v$_13554_out0 = v$A_11252_out0[11:11];
assign v$G3_206_out0 = ((v$_3282_out0 && !v$SUB_4616_out0) || (!v$_3282_out0) && v$SUB_4616_out0);
assign v$G3_208_out0 = ((v$_3284_out0 && !v$SUB_4618_out0) || (!v$_3284_out0) && v$SUB_4618_out0);
assign v$G8_549_out0 = v$_13385_out0 && v$_198_out0;
assign v$G8_551_out0 = v$_13387_out0 && v$_199_out0;
assign v$G14_616_out0 = v$_4712_out0 && v$_10538_out0;
assign v$G14_618_out0 = v$_4714_out0 && v$_10539_out0;
assign v$G13_643_out0 = v$_2876_out0 && v$_11212_out0;
assign v$G13_645_out0 = v$_2878_out0 && v$_11213_out0;
assign v$G8_1215_out0 = ((v$_8827_out0 && !v$SUB_4616_out0) || (!v$_8827_out0) && v$SUB_4616_out0);
assign v$G8_1217_out0 = ((v$_8829_out0 && !v$SUB_4618_out0) || (!v$_8829_out0) && v$SUB_4618_out0);
assign v$S_1240_out0 = v$S_8909_out0;
assign v$S_1464_out0 = v$S_9373_out0;
assign v$G2_1810_out0 = v$_13513_out0 && v$_13251_out0;
assign v$G2_1812_out0 = v$_13515_out0 && v$_13252_out0;
assign v$G15_1814_out0 = ((v$_3119_out0 && !v$SUB_4616_out0) || (!v$_3119_out0) && v$SUB_4616_out0);
assign v$G15_1816_out0 = ((v$_3121_out0 && !v$SUB_4618_out0) || (!v$_3121_out0) && v$SUB_4618_out0);
assign v$G1_1880_out0 = v$_1894_out0 && v$_7070_out0;
assign v$G1_1882_out0 = v$_1896_out0 && v$_7071_out0;
assign v$G10_2641_out0 = v$_13628_out0 && v$_1904_out0;
assign v$G10_2643_out0 = v$_13630_out0 && v$_1905_out0;
assign v$G4_2768_out0 = v$_2880_out0 && v$_4610_out0;
assign v$G4_2770_out0 = v$_2882_out0 && v$_4611_out0;
assign v$G7_2779_out0 = ((v$_2418_out0 && !v$SUB_4616_out0) || (!v$_2418_out0) && v$SUB_4616_out0);
assign v$G7_2781_out0 = ((v$_2420_out0 && !v$SUB_4618_out0) || (!v$_2420_out0) && v$SUB_4618_out0);
assign v$G5_2784_out0 = v$_1_out0 && v$_4812_out0;
assign v$G5_2786_out0 = v$_3_out0 && v$_4813_out0;
assign v$G9_2896_out0 = v$_3248_out0 && v$_13392_out0;
assign v$G9_2898_out0 = v$_3250_out0 && v$_13393_out0;
assign v$G11_2938_out0 = v$_4598_out0 && v$_2943_out0;
assign v$G11_2940_out0 = v$_4600_out0 && v$_2944_out0;
assign v$G12_3345_out0 = ((v$_13552_out0 && !v$SUB_4616_out0) || (!v$_13552_out0) && v$SUB_4616_out0);
assign v$G12_3347_out0 = ((v$_13554_out0 && !v$SUB_4618_out0) || (!v$_13554_out0) && v$SUB_4618_out0);
assign v$G1_4016_out0 = v$CARRY_4908_out0 || v$CARRY_4907_out0;
assign v$G1_4240_out0 = v$CARRY_5372_out0 || v$CARRY_5371_out0;
assign v$G14_4533_out0 = ((v$_2093_out0 && !v$SUB_4616_out0) || (!v$_2093_out0) && v$SUB_4616_out0);
assign v$G14_4535_out0 = ((v$_2095_out0 && !v$SUB_4618_out0) || (!v$_2095_out0) && v$SUB_4618_out0);
assign v$G15_4655_out0 = v$_8849_out0 && v$_4814_out0;
assign v$G15_4657_out0 = v$_8851_out0 && v$_4815_out0;
assign v$G13_4705_out0 = ((v$_10777_out0 && !v$SUB_4616_out0) || (!v$_10777_out0) && v$SUB_4616_out0);
assign v$G13_4707_out0 = ((v$_10779_out0 && !v$SUB_4618_out0) || (!v$_10779_out0) && v$SUB_4618_out0);
assign v$G2_7025_out0 = ((v$_10385_out0 && !v$SUB_4616_out0) || (!v$_10385_out0) && v$SUB_4616_out0);
assign v$G2_7027_out0 = ((v$_10387_out0 && !v$SUB_4618_out0) || (!v$_10387_out0) && v$SUB_4618_out0);
assign v$G3_7088_out0 = v$_2151_out0 && v$_2462_out0;
assign v$G3_7090_out0 = v$_2153_out0 && v$_2463_out0;
assign v$G7_8656_out0 = v$_11150_out0 && v$_4833_out0;
assign v$G7_8658_out0 = v$_11152_out0 && v$_4834_out0;
assign v$G6_8835_out0 = v$_1693_out0 && v$_1722_out0;
assign v$G6_8837_out0 = v$_1695_out0 && v$_1723_out0;
assign v$G5_10568_out0 = ((v$_10695_out0 && !v$SUB_4616_out0) || (!v$_10695_out0) && v$SUB_4616_out0);
assign v$G5_10570_out0 = ((v$_10697_out0 && !v$SUB_4618_out0) || (!v$_10697_out0) && v$SUB_4618_out0);
assign v$G12_10689_out0 = v$_1748_out0 && v$_3237_out0;
assign v$G12_10691_out0 = v$_1750_out0 && v$_3238_out0;
assign v$G16_10907_out0 = v$_2761_out0 && v$_8831_out0;
assign v$G16_10909_out0 = v$_2763_out0 && v$_8832_out0;
assign v$G4_10997_out0 = ((v$_77_out0 && !v$SUB_4616_out0) || (!v$_77_out0) && v$SUB_4616_out0);
assign v$G4_10999_out0 = ((v$_79_out0 && !v$SUB_4618_out0) || (!v$_79_out0) && v$SUB_4618_out0);
assign v$G16_11034_out0 = ((v$_192_out0 && !v$SUB_4616_out0) || (!v$_192_out0) && v$SUB_4616_out0);
assign v$G16_11036_out0 = ((v$_194_out0 && !v$SUB_4618_out0) || (!v$_194_out0) && v$SUB_4618_out0);
assign v$G10_13215_out0 = ((v$_329_out0 && !v$SUB_4616_out0) || (!v$_329_out0) && v$SUB_4616_out0);
assign v$G10_13217_out0 = ((v$_331_out0 && !v$SUB_4618_out0) || (!v$_331_out0) && v$SUB_4618_out0);
assign v$G9_13285_out0 = ((v$_8748_out0 && !v$SUB_4616_out0) || (!v$_8748_out0) && v$SUB_4616_out0);
assign v$G9_13287_out0 = ((v$_8750_out0 && !v$SUB_4618_out0) || (!v$_8750_out0) && v$SUB_4618_out0);
assign v$G11_13342_out0 = ((v$_10862_out0 && !v$SUB_4616_out0) || (!v$_10862_out0) && v$SUB_4616_out0);
assign v$G11_13344_out0 = ((v$_10864_out0 && !v$SUB_4618_out0) || (!v$_10864_out0) && v$SUB_4618_out0);
assign v$G6_13637_out0 = ((v$_10377_out0 && !v$SUB_4616_out0) || (!v$_10377_out0) && v$SUB_4616_out0);
assign v$G6_13639_out0 = ((v$_10379_out0 && !v$SUB_4618_out0) || (!v$_10379_out0) && v$SUB_4618_out0);
assign v$G1_13757_out0 = ((v$_321_out0 && !v$SUB_4616_out0) || (!v$_321_out0) && v$SUB_4616_out0);
assign v$G1_13759_out0 = ((v$_323_out0 && !v$SUB_4618_out0) || (!v$_323_out0) && v$SUB_4618_out0);
assign v$_387_out0 = { v$G5_2784_out0,v$G6_8835_out0 };
assign v$_389_out0 = { v$G5_2786_out0,v$G6_8837_out0 };
assign v$_400_out0 = { v$G9_2896_out0,v$G10_2641_out0 };
assign v$_402_out0 = { v$G9_2898_out0,v$G10_2643_out0 };
assign v$COUT_708_out0 = v$G1_4016_out0;
assign v$COUT_932_out0 = v$G1_4240_out0;
assign v$_1951_out0 = { v$G1_13757_out0,v$G2_7025_out0 };
assign v$_1953_out0 = { v$G1_13759_out0,v$G2_7027_out0 };
assign v$_2946_out0 = { v$G15_4655_out0,v$G16_10907_out0 };
assign v$_2948_out0 = { v$G15_4657_out0,v$G16_10909_out0 };
assign v$_3216_out0 = { v$G1_1880_out0,v$G2_1810_out0 };
assign v$_3218_out0 = { v$G1_1882_out0,v$G2_1812_out0 };
assign v$_3279_out0 = { v$G3_7088_out0,v$G4_2768_out0 };
assign v$_3281_out0 = { v$G3_7090_out0,v$G4_2770_out0 };
assign v$_5803_out0 = { v$_6927_out0,v$S_1240_out0 };
assign v$_5818_out0 = { v$_6942_out0,v$S_1464_out0 };
assign v$_7136_out0 = { v$G13_643_out0,v$G14_616_out0 };
assign v$_7138_out0 = { v$G13_645_out0,v$G14_618_out0 };
assign v$_13262_out0 = { v$G11_2938_out0,v$G12_10689_out0 };
assign v$_13264_out0 = { v$G11_2940_out0,v$G12_10691_out0 };
assign v$_13771_out0 = { v$G7_8656_out0,v$G8_549_out0 };
assign v$_13773_out0 = { v$G7_8658_out0,v$G8_551_out0 };
assign v$_114_out0 = { v$_387_out0,v$_13771_out0 };
assign v$_116_out0 = { v$_389_out0,v$_13773_out0 };
assign v$_450_out0 = { v$_7136_out0,v$_2946_out0 };
assign v$_452_out0 = { v$_7138_out0,v$_2948_out0 };
assign v$_2346_out0 = { v$_400_out0,v$_13262_out0 };
assign v$_2348_out0 = { v$_402_out0,v$_13264_out0 };
assign v$_9804_out0 = { v$_1951_out0,v$G3_206_out0 };
assign v$_9806_out0 = { v$_1953_out0,v$G3_208_out0 };
assign v$CIN_9834_out0 = v$COUT_708_out0;
assign v$CIN_10058_out0 = v$COUT_932_out0;
assign v$_10373_out0 = { v$_3216_out0,v$_3279_out0 };
assign v$_10375_out0 = { v$_3218_out0,v$_3281_out0 };
assign v$_2685_out0 = { v$_10373_out0,v$_114_out0 };
assign v$_2687_out0 = { v$_10375_out0,v$_116_out0 };
assign v$_4450_out0 = { v$_2346_out0,v$_450_out0 };
assign v$_4452_out0 = { v$_2348_out0,v$_452_out0 };
assign v$RD_5918_out0 = v$CIN_9834_out0;
assign v$RD_6382_out0 = v$CIN_10058_out0;
assign v$_8687_out0 = { v$_9804_out0,v$G4_10997_out0 };
assign v$_8689_out0 = { v$_9806_out0,v$G4_10999_out0 };
assign v$_1868_out0 = { v$_2685_out0,v$_4450_out0 };
assign v$_1870_out0 = { v$_2687_out0,v$_4452_out0 };
assign v$_3251_out0 = { v$_8687_out0,v$G5_10568_out0 };
assign v$_3253_out0 = { v$_8689_out0,v$G5_10570_out0 };
assign v$G1_7773_out0 = ((v$RD_5918_out0 && !v$RM_11358_out0) || (!v$RD_5918_out0) && v$RM_11358_out0);
assign v$G1_8237_out0 = ((v$RD_6382_out0 && !v$RM_11822_out0) || (!v$RD_6382_out0) && v$RM_11822_out0);
assign v$G2_12309_out0 = v$RD_5918_out0 && v$RM_11358_out0;
assign v$G2_12773_out0 = v$RD_6382_out0 && v$RM_11822_out0;
assign v$ANDOUT_631_out0 = v$_1868_out0;
assign v$ANDOUT_633_out0 = v$_1870_out0;
assign v$CARRY_4918_out0 = v$G2_12309_out0;
assign v$CARRY_5382_out0 = v$G2_12773_out0;
assign v$S_8919_out0 = v$G1_7773_out0;
assign v$S_9383_out0 = v$G1_8237_out0;
assign v$_10298_out0 = { v$_3251_out0,v$G6_13637_out0 };
assign v$_10300_out0 = { v$_3253_out0,v$G6_13639_out0 };
assign v$_119_out0 = { v$_10298_out0,v$G7_2779_out0 };
assign v$_121_out0 = { v$_10300_out0,v$G7_2781_out0 };
assign v$S_1245_out0 = v$S_8919_out0;
assign v$S_1469_out0 = v$S_9383_out0;
assign v$G1_4021_out0 = v$CARRY_4918_out0 || v$CARRY_4917_out0;
assign v$G1_4245_out0 = v$CARRY_5382_out0 || v$CARRY_5381_out0;
assign v$COUT_713_out0 = v$G1_4021_out0;
assign v$COUT_937_out0 = v$G1_4245_out0;
assign v$_2027_out0 = { v$_5803_out0,v$S_1245_out0 };
assign v$_2042_out0 = { v$_5818_out0,v$S_1469_out0 };
assign v$_13790_out0 = { v$_119_out0,v$G8_1215_out0 };
assign v$_13792_out0 = { v$_121_out0,v$G8_1217_out0 };
assign v$_464_out0 = { v$_13790_out0,v$G9_13285_out0 };
assign v$_466_out0 = { v$_13792_out0,v$G9_13287_out0 };
assign v$CIN_9823_out0 = v$COUT_713_out0;
assign v$CIN_10047_out0 = v$COUT_937_out0;
assign v$_422_out0 = { v$_464_out0,v$G10_13215_out0 };
assign v$_424_out0 = { v$_466_out0,v$G10_13217_out0 };
assign v$RD_5894_out0 = v$CIN_9823_out0;
assign v$RD_6358_out0 = v$CIN_10047_out0;
assign v$_2834_out0 = { v$_422_out0,v$G11_13342_out0 };
assign v$_2836_out0 = { v$_424_out0,v$G11_13344_out0 };
assign v$G1_7749_out0 = ((v$RD_5894_out0 && !v$RM_11334_out0) || (!v$RD_5894_out0) && v$RM_11334_out0);
assign v$G1_8213_out0 = ((v$RD_6358_out0 && !v$RM_11798_out0) || (!v$RD_6358_out0) && v$RM_11798_out0);
assign v$G2_12285_out0 = v$RD_5894_out0 && v$RM_11334_out0;
assign v$G2_12749_out0 = v$RD_6358_out0 && v$RM_11798_out0;
assign v$CARRY_4894_out0 = v$G2_12285_out0;
assign v$CARRY_5358_out0 = v$G2_12749_out0;
assign v$S_8895_out0 = v$G1_7749_out0;
assign v$S_9359_out0 = v$G1_8213_out0;
assign v$_11137_out0 = { v$_2834_out0,v$G12_3345_out0 };
assign v$_11139_out0 = { v$_2836_out0,v$G12_3347_out0 };
assign v$S_1234_out0 = v$S_8895_out0;
assign v$S_1458_out0 = v$S_9359_out0;
assign v$_3192_out0 = { v$_11137_out0,v$G13_4705_out0 };
assign v$_3194_out0 = { v$_11139_out0,v$G13_4707_out0 };
assign v$G1_4010_out0 = v$CARRY_4894_out0 || v$CARRY_4893_out0;
assign v$G1_4234_out0 = v$CARRY_5358_out0 || v$CARRY_5357_out0;
assign v$_173_out0 = { v$_3192_out0,v$G14_4533_out0 };
assign v$_175_out0 = { v$_3194_out0,v$G14_4535_out0 };
assign v$COUT_702_out0 = v$G1_4010_out0;
assign v$COUT_926_out0 = v$G1_4234_out0;
assign v$_2794_out0 = { v$_2027_out0,v$S_1234_out0 };
assign v$_2809_out0 = { v$_2042_out0,v$S_1458_out0 };
assign v$CIN_9827_out0 = v$COUT_702_out0;
assign v$CIN_10051_out0 = v$COUT_926_out0;
assign v$_10455_out0 = { v$_173_out0,v$G15_1814_out0 };
assign v$_10457_out0 = { v$_175_out0,v$G15_1816_out0 };
assign v$_1211_out0 = { v$_10455_out0,v$G16_11034_out0 };
assign v$_1213_out0 = { v$_10457_out0,v$G16_11036_out0 };
assign v$RD_5902_out0 = v$CIN_9827_out0;
assign v$RD_6366_out0 = v$CIN_10051_out0;
assign v$G1_7757_out0 = ((v$RD_5902_out0 && !v$RM_11342_out0) || (!v$RD_5902_out0) && v$RM_11342_out0);
assign v$G1_8221_out0 = ((v$RD_6366_out0 && !v$RM_11806_out0) || (!v$RD_6366_out0) && v$RM_11806_out0);
assign v$ADDER$IN_8744_out0 = v$_1211_out0;
assign v$ADDER$IN_8746_out0 = v$_1213_out0;
assign v$G2_12293_out0 = v$RD_5902_out0 && v$RM_11342_out0;
assign v$G2_12757_out0 = v$RD_6366_out0 && v$RM_11806_out0;
assign {v$A1_3855_out1,v$A1_3855_out0 } = v$OP1_2060_out0 + v$ADDER$IN_8744_out0 + v$G10_130_out0;
assign {v$A1_3856_out1,v$A1_3856_out0 } = v$OP1_2061_out0 + v$ADDER$IN_8746_out0 + v$G10_131_out0;
assign v$CARRY_4902_out0 = v$G2_12293_out0;
assign v$CARRY_5366_out0 = v$G2_12757_out0;
assign v$S_8903_out0 = v$G1_7757_out0;
assign v$S_9367_out0 = v$G1_8221_out0;
assign v$S_1238_out0 = v$S_8903_out0;
assign v$S_1462_out0 = v$S_9367_out0;
assign v$COUT_3895_out0 = v$A1_3855_out1;
assign v$COUT_3896_out0 = v$A1_3856_out1;
assign v$G1_4014_out0 = v$CARRY_4902_out0 || v$CARRY_4901_out0;
assign v$G1_4238_out0 = v$CARRY_5366_out0 || v$CARRY_5365_out0;
assign v$SUM1_13213_out0 = v$A1_3855_out0;
assign v$SUM1_13214_out0 = v$A1_3856_out0;
assign v$COUT_706_out0 = v$G1_4014_out0;
assign v$COUT_930_out0 = v$G1_4238_out0;
assign v$_1826_out0 = { v$_2794_out0,v$S_1238_out0 };
assign v$_1841_out0 = { v$_2809_out0,v$S_1462_out0 };
assign v$MUX3_2058_out0 = v$G7_169_out0 ? v$SUM1_13213_out0 : v$MUX5_2595_out0;
assign v$MUX3_2059_out0 = v$G7_170_out0 ? v$SUM1_13214_out0 : v$MUX5_2596_out0;
assign v$MUX2_1199_out0 = v$G9_411_out0 ? v$ANDOUT_631_out0 : v$MUX3_2058_out0;
assign v$MUX2_1200_out0 = v$G9_412_out0 ? v$ANDOUT_633_out0 : v$MUX3_2059_out0;
assign v$CIN_9824_out0 = v$COUT_706_out0;
assign v$CIN_10048_out0 = v$COUT_930_out0;
assign v$RD_5896_out0 = v$CIN_9824_out0;
assign v$RD_6360_out0 = v$CIN_10048_out0;
assign v$ALUOUT_10528_out0 = v$MUX2_1199_out0;
assign v$ALUOUT_10529_out0 = v$MUX2_1200_out0;
assign v$G1_7751_out0 = ((v$RD_5896_out0 && !v$RM_11336_out0) || (!v$RD_5896_out0) && v$RM_11336_out0);
assign v$G1_8215_out0 = ((v$RD_6360_out0 && !v$RM_11800_out0) || (!v$RD_6360_out0) && v$RM_11800_out0);
assign v$ALUOUT_8856_out0 = v$ALUOUT_10528_out0;
assign v$ALUOUT_8857_out0 = v$ALUOUT_10529_out0;
assign v$G2_12287_out0 = v$RD_5896_out0 && v$RM_11336_out0;
assign v$G2_12751_out0 = v$RD_6360_out0 && v$RM_11800_out0;
assign v$ALUOUT_4607_out0 = v$ALUOUT_8856_out0;
assign v$ALUOUT_4608_out0 = v$ALUOUT_8857_out0;
assign v$CARRY_4896_out0 = v$G2_12287_out0;
assign v$CARRY_5360_out0 = v$G2_12751_out0;
assign v$S_8897_out0 = v$G1_7751_out0;
assign v$S_9361_out0 = v$G1_8215_out0;
assign v$S_1235_out0 = v$S_8897_out0;
assign v$S_1459_out0 = v$S_9361_out0;
assign v$G1_4011_out0 = v$CARRY_4896_out0 || v$CARRY_4895_out0;
assign v$G1_4235_out0 = v$CARRY_5360_out0 || v$CARRY_5359_out0;
assign v$ALUOUT_11053_out0 = v$ALUOUT_4607_out0;
assign v$ALUOUT_11054_out0 = v$ALUOUT_4608_out0;
assign v$COUT_703_out0 = v$G1_4011_out0;
assign v$COUT_927_out0 = v$G1_4235_out0;
assign v$ALUOUT_4494_out0 = v$ALUOUT_11053_out0;
assign v$ALUOUT_4495_out0 = v$ALUOUT_11054_out0;
assign v$_4550_out0 = { v$_1826_out0,v$S_1235_out0 };
assign v$_4565_out0 = { v$_1841_out0,v$S_1459_out0 };
assign v$EQ3_11044_out0 = v$ALUOUT_4494_out0 == 16'h0;
assign v$EQ3_11045_out0 = v$ALUOUT_4495_out0 == 16'h0;
assign v$_11294_out0 = v$ALUOUT_4494_out0[14:0];
assign v$_11294_out1 = v$ALUOUT_4494_out0[15:1];
assign v$_11295_out0 = v$ALUOUT_4495_out0[14:0];
assign v$_11295_out1 = v$ALUOUT_4495_out0[15:1];
assign v$RM_11344_out0 = v$COUT_703_out0;
assign v$RM_11808_out0 = v$COUT_927_out0;
assign v$EQ_100_out0 = v$EQ3_11044_out0;
assign v$EQ_101_out0 = v$EQ3_11045_out0;
assign v$REST_162_out0 = v$_11294_out0;
assign v$REST_163_out0 = v$_11295_out0;
assign v$MI_2612_out0 = v$_11294_out1;
assign v$MI_2613_out0 = v$_11295_out1;
assign v$G1_7759_out0 = ((v$RD_5904_out0 && !v$RM_11344_out0) || (!v$RD_5904_out0) && v$RM_11344_out0);
assign v$G1_8223_out0 = ((v$RD_6368_out0 && !v$RM_11808_out0) || (!v$RD_6368_out0) && v$RM_11808_out0);
assign v$G2_12295_out0 = v$RD_5904_out0 && v$RM_11344_out0;
assign v$G2_12759_out0 = v$RD_6368_out0 && v$RM_11808_out0;
assign v$MI_560_out0 = v$MI_2612_out0;
assign v$MI_561_out0 = v$MI_2613_out0;
assign v$EQ_2591_out0 = v$EQ_100_out0;
assign v$EQ_2592_out0 = v$EQ_101_out0;
assign v$CARRY_4904_out0 = v$G2_12295_out0;
assign v$CARRY_5368_out0 = v$G2_12759_out0;
assign v$S_8905_out0 = v$G1_7759_out0;
assign v$S_9369_out0 = v$G1_8223_out0;
assign v$EQ_3821_out0 = v$EQ_2591_out0;
assign v$EQ_3822_out0 = v$EQ_2592_out0;
assign v$_10652_out0 = { v$_4550_out0,v$S_8905_out0 };
assign v$_10667_out0 = { v$_4565_out0,v$S_9369_out0 };
assign v$MI_10833_out0 = v$MI_560_out0;
assign v$MI_10834_out0 = v$MI_561_out0;
assign v$JMIN_2662_out0 = v$MI_10833_out0;
assign v$JMIN_2663_out0 = v$MI_10834_out0;
assign v$JEQZ_10514_out0 = v$EQ_3821_out0;
assign v$JEQZ_10515_out0 = v$EQ_3822_out0;
assign v$_10947_out0 = { v$_10652_out0,v$CARRY_4904_out0 };
assign v$_10962_out0 = { v$_10667_out0,v$CARRY_5368_out0 };
assign v$JMIN_1205_out0 = v$JMIN_2662_out0;
assign v$JMIN_1206_out0 = v$JMIN_2663_out0;
assign v$JEQZ_2981_out0 = v$JEQZ_10514_out0;
assign v$JEQZ_2982_out0 = v$JEQZ_10515_out0;
assign v$COUT_10917_out0 = v$_10947_out0;
assign v$COUT_10932_out0 = v$_10962_out0;
assign v$CIN_2357_out0 = v$COUT_10917_out0;
assign v$CIN_2372_out0 = v$COUT_10932_out0;
assign v$G4_4846_out0 = v$JEQZ_2981_out0 && v$JEQ_8806_out0;
assign v$G4_4847_out0 = v$JEQZ_2982_out0 && v$JEQ_8807_out0;
assign v$G5_10533_out0 = v$JMIN_1205_out0 && v$JMI_3212_out0;
assign v$G5_10534_out0 = v$JMIN_1206_out0 && v$JMI_3213_out0;
assign v$_470_out0 = v$CIN_2357_out0[8:8];
assign v$_485_out0 = v$CIN_2372_out0[8:8];
assign v$_1775_out0 = v$CIN_2357_out0[6:6];
assign v$_1790_out0 = v$CIN_2372_out0[6:6];
assign v$_2157_out0 = v$CIN_2357_out0[3:3];
assign v$_2172_out0 = v$CIN_2372_out0[3:3];
assign v$_2196_out0 = v$CIN_2357_out0[15:15];
assign v$_2210_out0 = v$CIN_2372_out0[15:15];
assign v$_2504_out0 = v$CIN_2357_out0[0:0];
assign v$_2519_out0 = v$CIN_2372_out0[0:0];
assign v$_3053_out0 = v$CIN_2357_out0[9:9];
assign v$_3068_out0 = v$CIN_2372_out0[9:9];
assign v$_3087_out0 = v$CIN_2357_out0[2:2];
assign v$_3102_out0 = v$CIN_2372_out0[2:2];
assign v$_3141_out0 = v$CIN_2357_out0[7:7];
assign v$_3156_out0 = v$CIN_2372_out0[7:7];
assign v$_3825_out0 = v$CIN_2357_out0[1:1];
assign v$_3840_out0 = v$CIN_2372_out0[1:1];
assign v$_3863_out0 = v$CIN_2357_out0[10:10];
assign v$_3878_out0 = v$CIN_2372_out0[10:10];
assign v$_6802_out0 = v$CIN_2357_out0[11:11];
assign v$_6817_out0 = v$CIN_2372_out0[11:11];
assign v$_7646_out0 = v$CIN_2357_out0[12:12];
assign v$_7661_out0 = v$CIN_2372_out0[12:12];
assign v$_8701_out0 = v$CIN_2357_out0[13:13];
assign v$_8716_out0 = v$CIN_2372_out0[13:13];
assign v$_8771_out0 = v$CIN_2357_out0[14:14];
assign v$_8786_out0 = v$CIN_2372_out0[14:14];
assign v$_10721_out0 = v$CIN_2357_out0[5:5];
assign v$_10736_out0 = v$CIN_2372_out0[5:5];
assign v$_13450_out0 = v$CIN_2357_out0[4:4];
assign v$_13465_out0 = v$CIN_2372_out0[4:4];
assign v$G2_13645_out0 = v$JMP_546_out0 || v$G5_10533_out0;
assign v$G2_13646_out0 = v$JMP_547_out0 || v$G5_10534_out0;
assign v$RM_3384_out0 = v$_7646_out0;
assign v$RM_3385_out0 = v$_8771_out0;
assign v$RM_3387_out0 = v$_10721_out0;
assign v$RM_3388_out0 = v$_13450_out0;
assign v$RM_3389_out0 = v$_8701_out0;
assign v$RM_3390_out0 = v$_3053_out0;
assign v$RM_3391_out0 = v$_3863_out0;
assign v$RM_3392_out0 = v$_3825_out0;
assign v$RM_3393_out0 = v$_2157_out0;
assign v$RM_3394_out0 = v$_1775_out0;
assign v$RM_3395_out0 = v$_3141_out0;
assign v$RM_3396_out0 = v$_6802_out0;
assign v$RM_3397_out0 = v$_470_out0;
assign v$RM_3398_out0 = v$_3087_out0;
assign v$RM_3608_out0 = v$_7661_out0;
assign v$RM_3609_out0 = v$_8786_out0;
assign v$RM_3611_out0 = v$_10736_out0;
assign v$RM_3612_out0 = v$_13465_out0;
assign v$RM_3613_out0 = v$_8716_out0;
assign v$RM_3614_out0 = v$_3068_out0;
assign v$RM_3615_out0 = v$_3878_out0;
assign v$RM_3616_out0 = v$_3840_out0;
assign v$RM_3617_out0 = v$_2172_out0;
assign v$RM_3618_out0 = v$_1790_out0;
assign v$RM_3619_out0 = v$_3156_out0;
assign v$RM_3620_out0 = v$_6817_out0;
assign v$RM_3621_out0 = v$_485_out0;
assign v$RM_3622_out0 = v$_3102_out0;
assign v$G3_3812_out0 = v$G2_13645_out0 || v$G4_4846_out0;
assign v$G3_3813_out0 = v$G2_13646_out0 || v$G4_4847_out0;
assign v$CIN_9839_out0 = v$_2196_out0;
assign v$CIN_10063_out0 = v$_2210_out0;
assign v$RM_11375_out0 = v$_2504_out0;
assign v$RM_11839_out0 = v$_2519_out0;
assign v$JUMP_2187_out0 = v$G3_3812_out0;
assign v$JUMP_2188_out0 = v$G3_3813_out0;
assign v$RD_5928_out0 = v$CIN_9839_out0;
assign v$RD_6392_out0 = v$CIN_10063_out0;
assign v$G1_7790_out0 = ((v$RD_5935_out0 && !v$RM_11375_out0) || (!v$RD_5935_out0) && v$RM_11375_out0);
assign v$G1_8254_out0 = ((v$RD_6399_out0 && !v$RM_11839_out0) || (!v$RD_6399_out0) && v$RM_11839_out0);
assign v$RM_11363_out0 = v$RM_3384_out0;
assign v$RM_11365_out0 = v$RM_3385_out0;
assign v$RM_11369_out0 = v$RM_3387_out0;
assign v$RM_11371_out0 = v$RM_3388_out0;
assign v$RM_11373_out0 = v$RM_3389_out0;
assign v$RM_11376_out0 = v$RM_3390_out0;
assign v$RM_11378_out0 = v$RM_3391_out0;
assign v$RM_11380_out0 = v$RM_3392_out0;
assign v$RM_11382_out0 = v$RM_3393_out0;
assign v$RM_11384_out0 = v$RM_3394_out0;
assign v$RM_11386_out0 = v$RM_3395_out0;
assign v$RM_11388_out0 = v$RM_3396_out0;
assign v$RM_11390_out0 = v$RM_3397_out0;
assign v$RM_11392_out0 = v$RM_3398_out0;
assign v$RM_11827_out0 = v$RM_3608_out0;
assign v$RM_11829_out0 = v$RM_3609_out0;
assign v$RM_11833_out0 = v$RM_3611_out0;
assign v$RM_11835_out0 = v$RM_3612_out0;
assign v$RM_11837_out0 = v$RM_3613_out0;
assign v$RM_11840_out0 = v$RM_3614_out0;
assign v$RM_11842_out0 = v$RM_3615_out0;
assign v$RM_11844_out0 = v$RM_3616_out0;
assign v$RM_11846_out0 = v$RM_3617_out0;
assign v$RM_11848_out0 = v$RM_3618_out0;
assign v$RM_11850_out0 = v$RM_3619_out0;
assign v$RM_11852_out0 = v$RM_3620_out0;
assign v$RM_11854_out0 = v$RM_3621_out0;
assign v$RM_11856_out0 = v$RM_3622_out0;
assign v$G2_12326_out0 = v$RD_5935_out0 && v$RM_11375_out0;
assign v$G2_12790_out0 = v$RD_6399_out0 && v$RM_11839_out0;
assign v$G14_1178_out0 = v$G15_1855_out0 && v$JUMP_2187_out0;
assign v$G14_1179_out0 = v$G15_1856_out0 && v$JUMP_2188_out0;
assign v$CARRY_4935_out0 = v$G2_12326_out0;
assign v$CARRY_5399_out0 = v$G2_12790_out0;
assign v$G1_7778_out0 = ((v$RD_5923_out0 && !v$RM_11363_out0) || (!v$RD_5923_out0) && v$RM_11363_out0);
assign v$G1_7780_out0 = ((v$RD_5925_out0 && !v$RM_11365_out0) || (!v$RD_5925_out0) && v$RM_11365_out0);
assign v$G1_7784_out0 = ((v$RD_5929_out0 && !v$RM_11369_out0) || (!v$RD_5929_out0) && v$RM_11369_out0);
assign v$G1_7786_out0 = ((v$RD_5931_out0 && !v$RM_11371_out0) || (!v$RD_5931_out0) && v$RM_11371_out0);
assign v$G1_7788_out0 = ((v$RD_5933_out0 && !v$RM_11373_out0) || (!v$RD_5933_out0) && v$RM_11373_out0);
assign v$G1_7791_out0 = ((v$RD_5936_out0 && !v$RM_11376_out0) || (!v$RD_5936_out0) && v$RM_11376_out0);
assign v$G1_7793_out0 = ((v$RD_5938_out0 && !v$RM_11378_out0) || (!v$RD_5938_out0) && v$RM_11378_out0);
assign v$G1_7795_out0 = ((v$RD_5940_out0 && !v$RM_11380_out0) || (!v$RD_5940_out0) && v$RM_11380_out0);
assign v$G1_7797_out0 = ((v$RD_5942_out0 && !v$RM_11382_out0) || (!v$RD_5942_out0) && v$RM_11382_out0);
assign v$G1_7799_out0 = ((v$RD_5944_out0 && !v$RM_11384_out0) || (!v$RD_5944_out0) && v$RM_11384_out0);
assign v$G1_7801_out0 = ((v$RD_5946_out0 && !v$RM_11386_out0) || (!v$RD_5946_out0) && v$RM_11386_out0);
assign v$G1_7803_out0 = ((v$RD_5948_out0 && !v$RM_11388_out0) || (!v$RD_5948_out0) && v$RM_11388_out0);
assign v$G1_7805_out0 = ((v$RD_5950_out0 && !v$RM_11390_out0) || (!v$RD_5950_out0) && v$RM_11390_out0);
assign v$G1_7807_out0 = ((v$RD_5952_out0 && !v$RM_11392_out0) || (!v$RD_5952_out0) && v$RM_11392_out0);
assign v$G1_8242_out0 = ((v$RD_6387_out0 && !v$RM_11827_out0) || (!v$RD_6387_out0) && v$RM_11827_out0);
assign v$G1_8244_out0 = ((v$RD_6389_out0 && !v$RM_11829_out0) || (!v$RD_6389_out0) && v$RM_11829_out0);
assign v$G1_8248_out0 = ((v$RD_6393_out0 && !v$RM_11833_out0) || (!v$RD_6393_out0) && v$RM_11833_out0);
assign v$G1_8250_out0 = ((v$RD_6395_out0 && !v$RM_11835_out0) || (!v$RD_6395_out0) && v$RM_11835_out0);
assign v$G1_8252_out0 = ((v$RD_6397_out0 && !v$RM_11837_out0) || (!v$RD_6397_out0) && v$RM_11837_out0);
assign v$G1_8255_out0 = ((v$RD_6400_out0 && !v$RM_11840_out0) || (!v$RD_6400_out0) && v$RM_11840_out0);
assign v$G1_8257_out0 = ((v$RD_6402_out0 && !v$RM_11842_out0) || (!v$RD_6402_out0) && v$RM_11842_out0);
assign v$G1_8259_out0 = ((v$RD_6404_out0 && !v$RM_11844_out0) || (!v$RD_6404_out0) && v$RM_11844_out0);
assign v$G1_8261_out0 = ((v$RD_6406_out0 && !v$RM_11846_out0) || (!v$RD_6406_out0) && v$RM_11846_out0);
assign v$G1_8263_out0 = ((v$RD_6408_out0 && !v$RM_11848_out0) || (!v$RD_6408_out0) && v$RM_11848_out0);
assign v$G1_8265_out0 = ((v$RD_6410_out0 && !v$RM_11850_out0) || (!v$RD_6410_out0) && v$RM_11850_out0);
assign v$G1_8267_out0 = ((v$RD_6412_out0 && !v$RM_11852_out0) || (!v$RD_6412_out0) && v$RM_11852_out0);
assign v$G1_8269_out0 = ((v$RD_6414_out0 && !v$RM_11854_out0) || (!v$RD_6414_out0) && v$RM_11854_out0);
assign v$G1_8271_out0 = ((v$RD_6416_out0 && !v$RM_11856_out0) || (!v$RD_6416_out0) && v$RM_11856_out0);
assign v$S_8936_out0 = v$G1_7790_out0;
assign v$S_9400_out0 = v$G1_8254_out0;
assign v$G2_12314_out0 = v$RD_5923_out0 && v$RM_11363_out0;
assign v$G2_12316_out0 = v$RD_5925_out0 && v$RM_11365_out0;
assign v$G2_12320_out0 = v$RD_5929_out0 && v$RM_11369_out0;
assign v$G2_12322_out0 = v$RD_5931_out0 && v$RM_11371_out0;
assign v$G2_12324_out0 = v$RD_5933_out0 && v$RM_11373_out0;
assign v$G2_12327_out0 = v$RD_5936_out0 && v$RM_11376_out0;
assign v$G2_12329_out0 = v$RD_5938_out0 && v$RM_11378_out0;
assign v$G2_12331_out0 = v$RD_5940_out0 && v$RM_11380_out0;
assign v$G2_12333_out0 = v$RD_5942_out0 && v$RM_11382_out0;
assign v$G2_12335_out0 = v$RD_5944_out0 && v$RM_11384_out0;
assign v$G2_12337_out0 = v$RD_5946_out0 && v$RM_11386_out0;
assign v$G2_12339_out0 = v$RD_5948_out0 && v$RM_11388_out0;
assign v$G2_12341_out0 = v$RD_5950_out0 && v$RM_11390_out0;
assign v$G2_12343_out0 = v$RD_5952_out0 && v$RM_11392_out0;
assign v$G2_12778_out0 = v$RD_6387_out0 && v$RM_11827_out0;
assign v$G2_12780_out0 = v$RD_6389_out0 && v$RM_11829_out0;
assign v$G2_12784_out0 = v$RD_6393_out0 && v$RM_11833_out0;
assign v$G2_12786_out0 = v$RD_6395_out0 && v$RM_11835_out0;
assign v$G2_12788_out0 = v$RD_6397_out0 && v$RM_11837_out0;
assign v$G2_12791_out0 = v$RD_6400_out0 && v$RM_11840_out0;
assign v$G2_12793_out0 = v$RD_6402_out0 && v$RM_11842_out0;
assign v$G2_12795_out0 = v$RD_6404_out0 && v$RM_11844_out0;
assign v$G2_12797_out0 = v$RD_6406_out0 && v$RM_11846_out0;
assign v$G2_12799_out0 = v$RD_6408_out0 && v$RM_11848_out0;
assign v$G2_12801_out0 = v$RD_6410_out0 && v$RM_11850_out0;
assign v$G2_12803_out0 = v$RD_6412_out0 && v$RM_11852_out0;
assign v$G2_12805_out0 = v$RD_6414_out0 && v$RM_11854_out0;
assign v$G2_12807_out0 = v$RD_6416_out0 && v$RM_11856_out0;
assign v$S_4667_out0 = v$S_8936_out0;
assign v$S_4682_out0 = v$S_9400_out0;
assign v$CARRY_4923_out0 = v$G2_12314_out0;
assign v$CARRY_4925_out0 = v$G2_12316_out0;
assign v$CARRY_4929_out0 = v$G2_12320_out0;
assign v$CARRY_4931_out0 = v$G2_12322_out0;
assign v$CARRY_4933_out0 = v$G2_12324_out0;
assign v$CARRY_4936_out0 = v$G2_12327_out0;
assign v$CARRY_4938_out0 = v$G2_12329_out0;
assign v$CARRY_4940_out0 = v$G2_12331_out0;
assign v$CARRY_4942_out0 = v$G2_12333_out0;
assign v$CARRY_4944_out0 = v$G2_12335_out0;
assign v$CARRY_4946_out0 = v$G2_12337_out0;
assign v$CARRY_4948_out0 = v$G2_12339_out0;
assign v$CARRY_4950_out0 = v$G2_12341_out0;
assign v$CARRY_4952_out0 = v$G2_12343_out0;
assign v$CARRY_5387_out0 = v$G2_12778_out0;
assign v$CARRY_5389_out0 = v$G2_12780_out0;
assign v$CARRY_5393_out0 = v$G2_12784_out0;
assign v$CARRY_5395_out0 = v$G2_12786_out0;
assign v$CARRY_5397_out0 = v$G2_12788_out0;
assign v$CARRY_5400_out0 = v$G2_12791_out0;
assign v$CARRY_5402_out0 = v$G2_12793_out0;
assign v$CARRY_5404_out0 = v$G2_12795_out0;
assign v$CARRY_5406_out0 = v$G2_12797_out0;
assign v$CARRY_5408_out0 = v$G2_12799_out0;
assign v$CARRY_5410_out0 = v$G2_12801_out0;
assign v$CARRY_5412_out0 = v$G2_12803_out0;
assign v$CARRY_5414_out0 = v$G2_12805_out0;
assign v$CARRY_5416_out0 = v$G2_12807_out0;
assign v$S_8924_out0 = v$G1_7778_out0;
assign v$S_8926_out0 = v$G1_7780_out0;
assign v$S_8930_out0 = v$G1_7784_out0;
assign v$S_8932_out0 = v$G1_7786_out0;
assign v$S_8934_out0 = v$G1_7788_out0;
assign v$S_8937_out0 = v$G1_7791_out0;
assign v$S_8939_out0 = v$G1_7793_out0;
assign v$S_8941_out0 = v$G1_7795_out0;
assign v$S_8943_out0 = v$G1_7797_out0;
assign v$S_8945_out0 = v$G1_7799_out0;
assign v$S_8947_out0 = v$G1_7801_out0;
assign v$S_8949_out0 = v$G1_7803_out0;
assign v$S_8951_out0 = v$G1_7805_out0;
assign v$S_8953_out0 = v$G1_7807_out0;
assign v$S_9388_out0 = v$G1_8242_out0;
assign v$S_9390_out0 = v$G1_8244_out0;
assign v$S_9394_out0 = v$G1_8248_out0;
assign v$S_9396_out0 = v$G1_8250_out0;
assign v$S_9398_out0 = v$G1_8252_out0;
assign v$S_9401_out0 = v$G1_8255_out0;
assign v$S_9403_out0 = v$G1_8257_out0;
assign v$S_9405_out0 = v$G1_8259_out0;
assign v$S_9407_out0 = v$G1_8261_out0;
assign v$S_9409_out0 = v$G1_8263_out0;
assign v$S_9411_out0 = v$G1_8265_out0;
assign v$S_9413_out0 = v$G1_8267_out0;
assign v$S_9415_out0 = v$G1_8269_out0;
assign v$S_9417_out0 = v$G1_8271_out0;
assign v$CIN_9845_out0 = v$CARRY_4935_out0;
assign v$CIN_10069_out0 = v$CARRY_5399_out0;
assign v$MUX1_10773_out0 = v$G14_1178_out0 ? v$JUMPADRESS_4745_out0 : v$REG1_432_out0;
assign v$MUX1_10774_out0 = v$G14_1179_out0 ? v$JUMPADRESS_4746_out0 : v$REG1_433_out0;
assign v$_1716_out0 = { v$_3223_out0,v$S_4667_out0 };
assign v$_1717_out0 = { v$_3224_out0,v$S_4682_out0 };
assign v$RD_5941_out0 = v$CIN_9845_out0;
assign v$RD_6405_out0 = v$CIN_10069_out0;
assign {v$A1_7019_out1,v$A1_7019_out0 } = v$MUX1_10773_out0 + v$ADDER$IN_10995_out0 + v$G22_1899_out0;
assign {v$A1_7020_out1,v$A1_7020_out0 } = v$MUX1_10774_out0 + v$ADDER$IN_10996_out0 + v$G22_1900_out0;
assign v$RM_11364_out0 = v$S_8924_out0;
assign v$RM_11366_out0 = v$S_8926_out0;
assign v$RM_11370_out0 = v$S_8930_out0;
assign v$RM_11372_out0 = v$S_8932_out0;
assign v$RM_11374_out0 = v$S_8934_out0;
assign v$RM_11377_out0 = v$S_8937_out0;
assign v$RM_11379_out0 = v$S_8939_out0;
assign v$RM_11381_out0 = v$S_8941_out0;
assign v$RM_11383_out0 = v$S_8943_out0;
assign v$RM_11385_out0 = v$S_8945_out0;
assign v$RM_11387_out0 = v$S_8947_out0;
assign v$RM_11389_out0 = v$S_8949_out0;
assign v$RM_11391_out0 = v$S_8951_out0;
assign v$RM_11393_out0 = v$S_8953_out0;
assign v$RM_11828_out0 = v$S_9388_out0;
assign v$RM_11830_out0 = v$S_9390_out0;
assign v$RM_11834_out0 = v$S_9394_out0;
assign v$RM_11836_out0 = v$S_9396_out0;
assign v$RM_11838_out0 = v$S_9398_out0;
assign v$RM_11841_out0 = v$S_9401_out0;
assign v$RM_11843_out0 = v$S_9403_out0;
assign v$RM_11845_out0 = v$S_9405_out0;
assign v$RM_11847_out0 = v$S_9407_out0;
assign v$RM_11849_out0 = v$S_9409_out0;
assign v$RM_11851_out0 = v$S_9411_out0;
assign v$RM_11853_out0 = v$S_9413_out0;
assign v$RM_11855_out0 = v$S_9415_out0;
assign v$RM_11857_out0 = v$S_9417_out0;
assign v$COUT_70_out0 = v$A1_7019_out1;
assign v$COUT_71_out0 = v$A1_7020_out1;
assign v$G1_7796_out0 = ((v$RD_5941_out0 && !v$RM_11381_out0) || (!v$RD_5941_out0) && v$RM_11381_out0);
assign v$G1_8260_out0 = ((v$RD_6405_out0 && !v$RM_11845_out0) || (!v$RD_6405_out0) && v$RM_11845_out0);
assign v$MUX3_10330_out0 = v$STP_11240_out0 ? v$A1_7019_out0 : v$MUX1_10773_out0;
assign v$MUX3_10331_out0 = v$STP_11241_out0 ? v$A1_7020_out0 : v$MUX1_10774_out0;
assign v$MUX5_10845_out0 = v$STORE$WEN_4544_out0 ? v$REG1_432_out0 : v$A1_7019_out0;
assign v$MUX5_10846_out0 = v$STORE$WEN_4545_out0 ? v$REG1_433_out0 : v$A1_7020_out0;
assign v$G2_12332_out0 = v$RD_5941_out0 && v$RM_11381_out0;
assign v$G2_12796_out0 = v$RD_6405_out0 && v$RM_11845_out0;
assign v$MUX4_2658_out0 = v$BYTE$READY_2852_out0 ? v$C1_2426_out0 : v$MUX5_10845_out0;
assign v$MUX4_2659_out0 = v$BYTE$READY_2853_out0 ? v$C1_2427_out0 : v$MUX5_10846_out0;
assign v$CARRY_4941_out0 = v$G2_12332_out0;
assign v$CARRY_5405_out0 = v$G2_12796_out0;
assign v$PC$COUNTER$NEXT_7064_out0 = v$MUX3_10330_out0;
assign v$PC$COUNTER$NEXT_7065_out0 = v$MUX3_10331_out0;
assign v$S_8942_out0 = v$G1_7796_out0;
assign v$S_9406_out0 = v$G1_8260_out0;
assign v$PC$COUNTER_25_out0 = v$PC$COUNTER$NEXT_7064_out0;
assign v$PC$COUNTER_26_out0 = v$PC$COUNTER$NEXT_7065_out0;
assign v$REGISTER_216_out0 = v$MUX4_2658_out0;
assign v$REGISTER_217_out0 = v$MUX4_2659_out0;
assign v$S_1256_out0 = v$S_8942_out0;
assign v$S_1480_out0 = v$S_9406_out0;
assign v$G1_4032_out0 = v$CARRY_4941_out0 || v$CARRY_4940_out0;
assign v$G1_4256_out0 = v$CARRY_5405_out0 || v$CARRY_5404_out0;
assign v$COUT_724_out0 = v$G1_4032_out0;
assign v$COUT_948_out0 = v$G1_4256_out0;
assign v$MUX3_3225_out0 = v$BYTE$READY_7021_out0 ? v$C2_10761_out0 : v$PC$COUNTER_25_out0;
assign v$MUX3_3226_out0 = v$BYTE$READY_7022_out0 ? v$C2_10762_out0 : v$PC$COUNTER_26_out0;
assign v$_8697_out0 = { v$PC$COUNTER_25_out0,v$C1_2005_out0 };
assign v$_8698_out0 = { v$PC$COUNTER_26_out0,v$C1_2006_out0 };
assign v$REGISTER_13346_out0 = v$REGISTER_216_out0;
assign v$REGISTER_13347_out0 = v$REGISTER_217_out0;
assign v$REGISTER4_1705_out0 = v$REGISTER_13346_out0;
assign v$REGISTER4_1706_out0 = v$REGISTER_13347_out0;
assign v$MUX2_3202_out0 = v$BYTE$READY_7021_out0 ? v$_8697_out0 : v$RAM$IN_233_out0;
assign v$MUX2_3203_out0 = v$BYTE$READY_7022_out0 ? v$_8698_out0 : v$RAM$IN_234_out0;
assign v$CIN_9851_out0 = v$COUT_724_out0;
assign v$CIN_10075_out0 = v$COUT_948_out0;
assign v$NEXTADD_10526_out0 = v$MUX3_3225_out0;
assign v$NEXTADD_10527_out0 = v$MUX3_3226_out0;
assign v$NEXTADRESS_1803_out0 = v$NEXTADD_10526_out0;
assign v$NEXTADRESS_1804_out0 = v$NEXTADD_10527_out0;
assign v$REGISTER14_3201_out0 = v$REGISTER4_1706_out0;
assign v$RD_5953_out0 = v$CIN_9851_out0;
assign v$RD_6417_out0 = v$CIN_10075_out0;
assign v$REGISTER15_8833_out0 = v$REGISTER4_1705_out0;
assign v$DATA$IN_10552_out0 = v$MUX2_3202_out0;
assign v$DATA$IN_10553_out0 = v$MUX2_3203_out0;
assign v$DATA$RAM$IN_558_out0 = v$DATA$IN_10552_out0;
assign v$DATA$RAM$IN_559_out0 = v$DATA$IN_10553_out0;
assign v$NEXT$ADRESS_3243_out0 = v$NEXTADRESS_1803_out0;
assign v$NEXT$ADRESS_3244_out0 = v$NEXTADRESS_1804_out0;
assign v$G1_7808_out0 = ((v$RD_5953_out0 && !v$RM_11393_out0) || (!v$RD_5953_out0) && v$RM_11393_out0);
assign v$G1_8272_out0 = ((v$RD_6417_out0 && !v$RM_11857_out0) || (!v$RD_6417_out0) && v$RM_11857_out0);
assign v$G2_12344_out0 = v$RD_5953_out0 && v$RM_11393_out0;
assign v$G2_12808_out0 = v$RD_6417_out0 && v$RM_11857_out0;
assign v$DATA$RAM$IN0_284_out0 = v$DATA$RAM$IN_559_out0;
assign v$DATA$RAM$IN1_4779_out0 = v$DATA$RAM$IN_558_out0;
assign v$CARRY_4953_out0 = v$G2_12344_out0;
assign v$CARRY_5417_out0 = v$G2_12808_out0;
assign v$S_8954_out0 = v$G1_7808_out0;
assign v$S_9418_out0 = v$G1_8272_out0;
assign v$ADRESS$ins1_10617_out0 = v$NEXT$ADRESS_3243_out0;
assign v$ADRESS$ins0_11169_out0 = v$NEXT$ADRESS_3244_out0;
assign v$DATA1_603_out0 = v$DATA$RAM$IN1_4779_out0;
assign v$S_1262_out0 = v$S_8954_out0;
assign v$S_1486_out0 = v$S_9418_out0;
assign v$G1_4038_out0 = v$CARRY_4953_out0 || v$CARRY_4952_out0;
assign v$G1_4262_out0 = v$CARRY_5417_out0 || v$CARRY_5416_out0;
assign v$DATA0_4737_out0 = v$DATA$RAM$IN0_284_out0;
assign v$COUT_730_out0 = v$G1_4038_out0;
assign v$COUT_954_out0 = v$G1_4262_out0;
assign v$DATA1_1974_out0 = v$DATA1_603_out0;
assign v$_4784_out0 = { v$S_1256_out0,v$S_1262_out0 };
assign v$_4799_out0 = { v$S_1480_out0,v$S_1486_out0 };
assign v$DATA0_13293_out0 = v$DATA0_4737_out0;
assign v$MUX4_1698_out0 = v$TX$inst0_608_out0 ? v$DATA0_13293_out0 : v$DATA1_1974_out0;
assign v$CIN_9846_out0 = v$COUT_730_out0;
assign v$CIN_10070_out0 = v$COUT_954_out0;
assign v$MUX3_10787_out0 = v$MUX$ENABLE_2349_out0 ? v$DATA0_13293_out0 : v$DATA1_1974_out0;
assign v$DATA$to$transmit_4546_out0 = v$MUX4_1698_out0;
assign v$RD_5943_out0 = v$CIN_9846_out0;
assign v$RD_6407_out0 = v$CIN_10070_out0;
assign v$DATA_10445_out0 = v$MUX3_10787_out0;
assign v$DATA_2469_out0 = v$DATA_10445_out0;
assign v$REGISTER$OUTPUT_3268_out0 = v$DATA$to$transmit_4546_out0;
assign v$G1_7798_out0 = ((v$RD_5943_out0 && !v$RM_11383_out0) || (!v$RD_5943_out0) && v$RM_11383_out0);
assign v$G1_8262_out0 = ((v$RD_6407_out0 && !v$RM_11847_out0) || (!v$RD_6407_out0) && v$RM_11847_out0);
assign v$G2_12334_out0 = v$RD_5943_out0 && v$RM_11383_out0;
assign v$G2_12798_out0 = v$RD_6407_out0 && v$RM_11847_out0;
assign v$REGISTER$OUTPUT2_2398_out0 = v$REGISTER$OUTPUT_3268_out0;
assign v$CARRY_4943_out0 = v$G2_12334_out0;
assign v$CARRY_5407_out0 = v$G2_12798_out0;
assign v$S_8944_out0 = v$G1_7798_out0;
assign v$S_9408_out0 = v$G1_8262_out0;
assign v$S_1257_out0 = v$S_8944_out0;
assign v$S_1481_out0 = v$S_9408_out0;
assign v$split_3196_out0 = v$REGISTER$OUTPUT2_2398_out0[7:0];
assign v$split_3196_out1 = v$REGISTER$OUTPUT2_2398_out0[15:8];
assign v$G1_4033_out0 = v$CARRY_4943_out0 || v$CARRY_4942_out0;
assign v$G1_4257_out0 = v$CARRY_5407_out0 || v$CARRY_5406_out0;
assign v$COUT_725_out0 = v$G1_4033_out0;
assign v$COUT_949_out0 = v$G1_4257_out0;
assign v$_2554_out0 = { v$_4784_out0,v$S_1257_out0 };
assign v$_2569_out0 = { v$_4799_out0,v$S_1481_out0 };
assign v$MUX1_13260_out0 = v$BYTE$COMP$1_8743_out0 ? v$split_3196_out1 : v$split_3196_out0;
assign v$TRANSMISSION$DATA2_7014_out0 = v$MUX1_13260_out0;
assign v$CIN_9841_out0 = v$COUT_725_out0;
assign v$CIN_10065_out0 = v$COUT_949_out0;
assign v$REGISTER$TRANSMIT$DATA_12241_out0 = v$MUX1_13260_out0;
assign v$TRANSMIT$DATA_76_out0 = v$REGISTER$TRANSMIT$DATA_12241_out0;
assign v$RD_5932_out0 = v$CIN_9841_out0;
assign v$RD_6396_out0 = v$CIN_10065_out0;
assign v$TRANSIMISSION$DATA_10818_out0 = v$TRANSMISSION$DATA2_7014_out0;
assign v$SEL1_240_out0 = v$TRANSMIT$DATA_76_out0[6:6];
assign v$SEL1_1164_out0 = v$TRANSMIT$DATA_76_out0[2:2];
assign v$SEL1_1204_out0 = v$TRANSMIT$DATA_76_out0[4:4];
assign v$SEL1_2319_out0 = v$TRANSMIT$DATA_76_out0[0:0];
assign v$SEL1_2428_out0 = v$TRANSMIT$DATA_76_out0[5:5];
assign v$SEL1_4858_out0 = v$TRANSMIT$DATA_76_out0[3:3];
assign v$G1_7787_out0 = ((v$RD_5932_out0 && !v$RM_11372_out0) || (!v$RD_5932_out0) && v$RM_11372_out0);
assign v$G1_8251_out0 = ((v$RD_6396_out0 && !v$RM_11836_out0) || (!v$RD_6396_out0) && v$RM_11836_out0);
assign v$SEL1_10304_out0 = v$TRANSMIT$DATA_76_out0[1:1];
assign v$G2_12323_out0 = v$RD_5932_out0 && v$RM_11372_out0;
assign v$G2_12787_out0 = v$RD_6396_out0 && v$RM_11836_out0;
assign v$SEL1_13445_out0 = v$TRANSMIT$DATA_76_out0[7:7];
assign v$MUX1_2625_out0 = v$transmit$INSTRUCTION_2674_out0 ? v$SEL1_240_out0 : v$FF1_1955_out0;
assign v$MUX4_3219_out0 = v$transmit$INSTRUCTION_2674_out0 ? v$SEL1_4858_out0 : v$FF4_463_out0;
assign v$MUX2_4448_out0 = v$transmit$INSTRUCTION_2674_out0 ? v$SEL1_2428_out0 : v$FF2_2833_out0;
assign v$CARRY_4932_out0 = v$G2_12323_out0;
assign v$CARRY_5396_out0 = v$G2_12787_out0;
assign v$MUX3_7140_out0 = v$transmit$INSTRUCTION_2674_out0 ? v$SEL1_1204_out0 : v$FF3_11046_out0;
assign v$S_8933_out0 = v$G1_7787_out0;
assign v$S_9397_out0 = v$G1_8251_out0;
assign v$MUX7_10448_out0 = v$transmit$INSTRUCTION_2674_out0 ? v$SEL1_2319_out0 : v$FF7_4781_out0;
assign v$MUX6_10976_out0 = v$transmit$INSTRUCTION_2674_out0 ? v$SEL1_10304_out0 : v$FF6_112_out0;
assign v$MUX5_13348_out0 = v$transmit$INSTRUCTION_2674_out0 ? v$SEL1_1164_out0 : v$FF5_7100_out0;
assign v$S_1252_out0 = v$S_8933_out0;
assign v$S_1476_out0 = v$S_9397_out0;
assign v$G1_4028_out0 = v$CARRY_4932_out0 || v$CARRY_4931_out0;
assign v$G1_4252_out0 = v$CARRY_5396_out0 || v$CARRY_5395_out0;
assign v$COUT_720_out0 = v$G1_4028_out0;
assign v$COUT_944_out0 = v$G1_4252_out0;
assign v$_7034_out0 = { v$_2554_out0,v$S_1252_out0 };
assign v$_7049_out0 = { v$_2569_out0,v$S_1476_out0 };
assign v$CIN_9840_out0 = v$COUT_720_out0;
assign v$CIN_10064_out0 = v$COUT_944_out0;
assign v$RD_5930_out0 = v$CIN_9840_out0;
assign v$RD_6394_out0 = v$CIN_10064_out0;
assign v$G1_7785_out0 = ((v$RD_5930_out0 && !v$RM_11370_out0) || (!v$RD_5930_out0) && v$RM_11370_out0);
assign v$G1_8249_out0 = ((v$RD_6394_out0 && !v$RM_11834_out0) || (!v$RD_6394_out0) && v$RM_11834_out0);
assign v$G2_12321_out0 = v$RD_5930_out0 && v$RM_11370_out0;
assign v$G2_12785_out0 = v$RD_6394_out0 && v$RM_11834_out0;
assign v$CARRY_4930_out0 = v$G2_12321_out0;
assign v$CARRY_5394_out0 = v$G2_12785_out0;
assign v$S_8931_out0 = v$G1_7785_out0;
assign v$S_9395_out0 = v$G1_8249_out0;
assign v$S_1251_out0 = v$S_8931_out0;
assign v$S_1475_out0 = v$S_9395_out0;
assign v$G1_4027_out0 = v$CARRY_4930_out0 || v$CARRY_4929_out0;
assign v$G1_4251_out0 = v$CARRY_5394_out0 || v$CARRY_5393_out0;
assign v$COUT_719_out0 = v$G1_4027_out0;
assign v$COUT_943_out0 = v$G1_4251_out0;
assign v$_13520_out0 = { v$_7034_out0,v$S_1251_out0 };
assign v$_13535_out0 = { v$_7049_out0,v$S_1475_out0 };
assign v$CIN_9847_out0 = v$COUT_719_out0;
assign v$CIN_10071_out0 = v$COUT_943_out0;
assign v$RD_5945_out0 = v$CIN_9847_out0;
assign v$RD_6409_out0 = v$CIN_10071_out0;
assign v$G1_7800_out0 = ((v$RD_5945_out0 && !v$RM_11385_out0) || (!v$RD_5945_out0) && v$RM_11385_out0);
assign v$G1_8264_out0 = ((v$RD_6409_out0 && !v$RM_11849_out0) || (!v$RD_6409_out0) && v$RM_11849_out0);
assign v$G2_12336_out0 = v$RD_5945_out0 && v$RM_11385_out0;
assign v$G2_12800_out0 = v$RD_6409_out0 && v$RM_11849_out0;
assign v$CARRY_4945_out0 = v$G2_12336_out0;
assign v$CARRY_5409_out0 = v$G2_12800_out0;
assign v$S_8946_out0 = v$G1_7800_out0;
assign v$S_9410_out0 = v$G1_8264_out0;
assign v$S_1258_out0 = v$S_8946_out0;
assign v$S_1482_out0 = v$S_9410_out0;
assign v$G1_4034_out0 = v$CARRY_4945_out0 || v$CARRY_4944_out0;
assign v$G1_4258_out0 = v$CARRY_5409_out0 || v$CARRY_5408_out0;
assign v$COUT_726_out0 = v$G1_4034_out0;
assign v$COUT_950_out0 = v$G1_4258_out0;
assign v$_3313_out0 = { v$_13520_out0,v$S_1258_out0 };
assign v$_3328_out0 = { v$_13535_out0,v$S_1482_out0 };
assign v$CIN_9848_out0 = v$COUT_726_out0;
assign v$CIN_10072_out0 = v$COUT_950_out0;
assign v$RD_5947_out0 = v$CIN_9848_out0;
assign v$RD_6411_out0 = v$CIN_10072_out0;
assign v$G1_7802_out0 = ((v$RD_5947_out0 && !v$RM_11387_out0) || (!v$RD_5947_out0) && v$RM_11387_out0);
assign v$G1_8266_out0 = ((v$RD_6411_out0 && !v$RM_11851_out0) || (!v$RD_6411_out0) && v$RM_11851_out0);
assign v$G2_12338_out0 = v$RD_5947_out0 && v$RM_11387_out0;
assign v$G2_12802_out0 = v$RD_6411_out0 && v$RM_11851_out0;
assign v$CARRY_4947_out0 = v$G2_12338_out0;
assign v$CARRY_5411_out0 = v$G2_12802_out0;
assign v$S_8948_out0 = v$G1_7802_out0;
assign v$S_9412_out0 = v$G1_8266_out0;
assign v$S_1259_out0 = v$S_8948_out0;
assign v$S_1483_out0 = v$S_9412_out0;
assign v$G1_4035_out0 = v$CARRY_4947_out0 || v$CARRY_4946_out0;
assign v$G1_4259_out0 = v$CARRY_5411_out0 || v$CARRY_5410_out0;
assign v$COUT_727_out0 = v$G1_4035_out0;
assign v$COUT_951_out0 = v$G1_4259_out0;
assign v$_7149_out0 = { v$_3313_out0,v$S_1259_out0 };
assign v$_7164_out0 = { v$_3328_out0,v$S_1483_out0 };
assign v$CIN_9850_out0 = v$COUT_727_out0;
assign v$CIN_10074_out0 = v$COUT_951_out0;
assign v$RD_5951_out0 = v$CIN_9850_out0;
assign v$RD_6415_out0 = v$CIN_10074_out0;
assign v$G1_7806_out0 = ((v$RD_5951_out0 && !v$RM_11391_out0) || (!v$RD_5951_out0) && v$RM_11391_out0);
assign v$G1_8270_out0 = ((v$RD_6415_out0 && !v$RM_11855_out0) || (!v$RD_6415_out0) && v$RM_11855_out0);
assign v$G2_12342_out0 = v$RD_5951_out0 && v$RM_11391_out0;
assign v$G2_12806_out0 = v$RD_6415_out0 && v$RM_11855_out0;
assign v$CARRY_4951_out0 = v$G2_12342_out0;
assign v$CARRY_5415_out0 = v$G2_12806_out0;
assign v$S_8952_out0 = v$G1_7806_out0;
assign v$S_9416_out0 = v$G1_8270_out0;
assign v$S_1261_out0 = v$S_8952_out0;
assign v$S_1485_out0 = v$S_9416_out0;
assign v$G1_4037_out0 = v$CARRY_4951_out0 || v$CARRY_4950_out0;
assign v$G1_4261_out0 = v$CARRY_5415_out0 || v$CARRY_5414_out0;
assign v$COUT_729_out0 = v$G1_4037_out0;
assign v$COUT_953_out0 = v$G1_4261_out0;
assign v$_4751_out0 = { v$_7149_out0,v$S_1261_out0 };
assign v$_4766_out0 = { v$_7164_out0,v$S_1485_out0 };
assign v$CIN_9843_out0 = v$COUT_729_out0;
assign v$CIN_10067_out0 = v$COUT_953_out0;
assign v$RD_5937_out0 = v$CIN_9843_out0;
assign v$RD_6401_out0 = v$CIN_10067_out0;
assign v$G1_7792_out0 = ((v$RD_5937_out0 && !v$RM_11377_out0) || (!v$RD_5937_out0) && v$RM_11377_out0);
assign v$G1_8256_out0 = ((v$RD_6401_out0 && !v$RM_11841_out0) || (!v$RD_6401_out0) && v$RM_11841_out0);
assign v$G2_12328_out0 = v$RD_5937_out0 && v$RM_11377_out0;
assign v$G2_12792_out0 = v$RD_6401_out0 && v$RM_11841_out0;
assign v$CARRY_4937_out0 = v$G2_12328_out0;
assign v$CARRY_5401_out0 = v$G2_12792_out0;
assign v$S_8938_out0 = v$G1_7792_out0;
assign v$S_9402_out0 = v$G1_8256_out0;
assign v$S_1254_out0 = v$S_8938_out0;
assign v$S_1478_out0 = v$S_9402_out0;
assign v$G1_4030_out0 = v$CARRY_4937_out0 || v$CARRY_4936_out0;
assign v$G1_4254_out0 = v$CARRY_5401_out0 || v$CARRY_5400_out0;
assign v$COUT_722_out0 = v$G1_4030_out0;
assign v$COUT_946_out0 = v$G1_4254_out0;
assign v$_6928_out0 = { v$_4751_out0,v$S_1254_out0 };
assign v$_6943_out0 = { v$_4766_out0,v$S_1478_out0 };
assign v$CIN_9844_out0 = v$COUT_722_out0;
assign v$CIN_10068_out0 = v$COUT_946_out0;
assign v$RD_5939_out0 = v$CIN_9844_out0;
assign v$RD_6403_out0 = v$CIN_10068_out0;
assign v$G1_7794_out0 = ((v$RD_5939_out0 && !v$RM_11379_out0) || (!v$RD_5939_out0) && v$RM_11379_out0);
assign v$G1_8258_out0 = ((v$RD_6403_out0 && !v$RM_11843_out0) || (!v$RD_6403_out0) && v$RM_11843_out0);
assign v$G2_12330_out0 = v$RD_5939_out0 && v$RM_11379_out0;
assign v$G2_12794_out0 = v$RD_6403_out0 && v$RM_11843_out0;
assign v$CARRY_4939_out0 = v$G2_12330_out0;
assign v$CARRY_5403_out0 = v$G2_12794_out0;
assign v$S_8940_out0 = v$G1_7794_out0;
assign v$S_9404_out0 = v$G1_8258_out0;
assign v$S_1255_out0 = v$S_8940_out0;
assign v$S_1479_out0 = v$S_9404_out0;
assign v$G1_4031_out0 = v$CARRY_4939_out0 || v$CARRY_4938_out0;
assign v$G1_4255_out0 = v$CARRY_5403_out0 || v$CARRY_5402_out0;
assign v$COUT_723_out0 = v$G1_4031_out0;
assign v$COUT_947_out0 = v$G1_4255_out0;
assign v$_5804_out0 = { v$_6928_out0,v$S_1255_out0 };
assign v$_5819_out0 = { v$_6943_out0,v$S_1479_out0 };
assign v$CIN_9849_out0 = v$COUT_723_out0;
assign v$CIN_10073_out0 = v$COUT_947_out0;
assign v$RD_5949_out0 = v$CIN_9849_out0;
assign v$RD_6413_out0 = v$CIN_10073_out0;
assign v$G1_7804_out0 = ((v$RD_5949_out0 && !v$RM_11389_out0) || (!v$RD_5949_out0) && v$RM_11389_out0);
assign v$G1_8268_out0 = ((v$RD_6413_out0 && !v$RM_11853_out0) || (!v$RD_6413_out0) && v$RM_11853_out0);
assign v$G2_12340_out0 = v$RD_5949_out0 && v$RM_11389_out0;
assign v$G2_12804_out0 = v$RD_6413_out0 && v$RM_11853_out0;
assign v$CARRY_4949_out0 = v$G2_12340_out0;
assign v$CARRY_5413_out0 = v$G2_12804_out0;
assign v$S_8950_out0 = v$G1_7804_out0;
assign v$S_9414_out0 = v$G1_8268_out0;
assign v$S_1260_out0 = v$S_8950_out0;
assign v$S_1484_out0 = v$S_9414_out0;
assign v$G1_4036_out0 = v$CARRY_4949_out0 || v$CARRY_4948_out0;
assign v$G1_4260_out0 = v$CARRY_5413_out0 || v$CARRY_5412_out0;
assign v$COUT_728_out0 = v$G1_4036_out0;
assign v$COUT_952_out0 = v$G1_4260_out0;
assign v$_2028_out0 = { v$_5804_out0,v$S_1260_out0 };
assign v$_2043_out0 = { v$_5819_out0,v$S_1484_out0 };
assign v$CIN_9837_out0 = v$COUT_728_out0;
assign v$CIN_10061_out0 = v$COUT_952_out0;
assign v$RD_5924_out0 = v$CIN_9837_out0;
assign v$RD_6388_out0 = v$CIN_10061_out0;
assign v$G1_7779_out0 = ((v$RD_5924_out0 && !v$RM_11364_out0) || (!v$RD_5924_out0) && v$RM_11364_out0);
assign v$G1_8243_out0 = ((v$RD_6388_out0 && !v$RM_11828_out0) || (!v$RD_6388_out0) && v$RM_11828_out0);
assign v$G2_12315_out0 = v$RD_5924_out0 && v$RM_11364_out0;
assign v$G2_12779_out0 = v$RD_6388_out0 && v$RM_11828_out0;
assign v$CARRY_4924_out0 = v$G2_12315_out0;
assign v$CARRY_5388_out0 = v$G2_12779_out0;
assign v$S_8925_out0 = v$G1_7779_out0;
assign v$S_9389_out0 = v$G1_8243_out0;
assign v$S_1248_out0 = v$S_8925_out0;
assign v$S_1472_out0 = v$S_9389_out0;
assign v$G1_4024_out0 = v$CARRY_4924_out0 || v$CARRY_4923_out0;
assign v$G1_4248_out0 = v$CARRY_5388_out0 || v$CARRY_5387_out0;
assign v$COUT_716_out0 = v$G1_4024_out0;
assign v$COUT_940_out0 = v$G1_4248_out0;
assign v$_2795_out0 = { v$_2028_out0,v$S_1248_out0 };
assign v$_2810_out0 = { v$_2043_out0,v$S_1472_out0 };
assign v$CIN_9842_out0 = v$COUT_716_out0;
assign v$CIN_10066_out0 = v$COUT_940_out0;
assign v$RD_5934_out0 = v$CIN_9842_out0;
assign v$RD_6398_out0 = v$CIN_10066_out0;
assign v$G1_7789_out0 = ((v$RD_5934_out0 && !v$RM_11374_out0) || (!v$RD_5934_out0) && v$RM_11374_out0);
assign v$G1_8253_out0 = ((v$RD_6398_out0 && !v$RM_11838_out0) || (!v$RD_6398_out0) && v$RM_11838_out0);
assign v$G2_12325_out0 = v$RD_5934_out0 && v$RM_11374_out0;
assign v$G2_12789_out0 = v$RD_6398_out0 && v$RM_11838_out0;
assign v$CARRY_4934_out0 = v$G2_12325_out0;
assign v$CARRY_5398_out0 = v$G2_12789_out0;
assign v$S_8935_out0 = v$G1_7789_out0;
assign v$S_9399_out0 = v$G1_8253_out0;
assign v$S_1253_out0 = v$S_8935_out0;
assign v$S_1477_out0 = v$S_9399_out0;
assign v$G1_4029_out0 = v$CARRY_4934_out0 || v$CARRY_4933_out0;
assign v$G1_4253_out0 = v$CARRY_5398_out0 || v$CARRY_5397_out0;
assign v$COUT_721_out0 = v$G1_4029_out0;
assign v$COUT_945_out0 = v$G1_4253_out0;
assign v$_1827_out0 = { v$_2795_out0,v$S_1253_out0 };
assign v$_1842_out0 = { v$_2810_out0,v$S_1477_out0 };
assign v$CIN_9838_out0 = v$COUT_721_out0;
assign v$CIN_10062_out0 = v$COUT_945_out0;
assign v$RD_5926_out0 = v$CIN_9838_out0;
assign v$RD_6390_out0 = v$CIN_10062_out0;
assign v$G1_7781_out0 = ((v$RD_5926_out0 && !v$RM_11366_out0) || (!v$RD_5926_out0) && v$RM_11366_out0);
assign v$G1_8245_out0 = ((v$RD_6390_out0 && !v$RM_11830_out0) || (!v$RD_6390_out0) && v$RM_11830_out0);
assign v$G2_12317_out0 = v$RD_5926_out0 && v$RM_11366_out0;
assign v$G2_12781_out0 = v$RD_6390_out0 && v$RM_11830_out0;
assign v$CARRY_4926_out0 = v$G2_12317_out0;
assign v$CARRY_5390_out0 = v$G2_12781_out0;
assign v$S_8927_out0 = v$G1_7781_out0;
assign v$S_9391_out0 = v$G1_8245_out0;
assign v$S_1249_out0 = v$S_8927_out0;
assign v$S_1473_out0 = v$S_9391_out0;
assign v$G1_4025_out0 = v$CARRY_4926_out0 || v$CARRY_4925_out0;
assign v$G1_4249_out0 = v$CARRY_5390_out0 || v$CARRY_5389_out0;
assign v$COUT_717_out0 = v$G1_4025_out0;
assign v$COUT_941_out0 = v$G1_4249_out0;
assign v$_4551_out0 = { v$_1827_out0,v$S_1249_out0 };
assign v$_4566_out0 = { v$_1842_out0,v$S_1473_out0 };
assign v$RM_3386_out0 = v$COUT_717_out0;
assign v$RM_3610_out0 = v$COUT_941_out0;
assign v$RM_11367_out0 = v$RM_3386_out0;
assign v$RM_11831_out0 = v$RM_3610_out0;
assign v$G1_7782_out0 = ((v$RD_5927_out0 && !v$RM_11367_out0) || (!v$RD_5927_out0) && v$RM_11367_out0);
assign v$G1_8246_out0 = ((v$RD_6391_out0 && !v$RM_11831_out0) || (!v$RD_6391_out0) && v$RM_11831_out0);
assign v$G2_12318_out0 = v$RD_5927_out0 && v$RM_11367_out0;
assign v$G2_12782_out0 = v$RD_6391_out0 && v$RM_11831_out0;
assign v$CARRY_4927_out0 = v$G2_12318_out0;
assign v$CARRY_5391_out0 = v$G2_12782_out0;
assign v$S_8928_out0 = v$G1_7782_out0;
assign v$S_9392_out0 = v$G1_8246_out0;
assign v$RM_11368_out0 = v$S_8928_out0;
assign v$RM_11832_out0 = v$S_9392_out0;
assign v$G1_7783_out0 = ((v$RD_5928_out0 && !v$RM_11368_out0) || (!v$RD_5928_out0) && v$RM_11368_out0);
assign v$G1_8247_out0 = ((v$RD_6392_out0 && !v$RM_11832_out0) || (!v$RD_6392_out0) && v$RM_11832_out0);
assign v$G2_12319_out0 = v$RD_5928_out0 && v$RM_11368_out0;
assign v$G2_12783_out0 = v$RD_6392_out0 && v$RM_11832_out0;
assign v$CARRY_4928_out0 = v$G2_12319_out0;
assign v$CARRY_5392_out0 = v$G2_12783_out0;
assign v$S_8929_out0 = v$G1_7783_out0;
assign v$S_9393_out0 = v$G1_8247_out0;
assign v$S_1250_out0 = v$S_8929_out0;
assign v$S_1474_out0 = v$S_9393_out0;
assign v$G1_4026_out0 = v$CARRY_4928_out0 || v$CARRY_4927_out0;
assign v$G1_4250_out0 = v$CARRY_5392_out0 || v$CARRY_5391_out0;
assign v$COUT_718_out0 = v$G1_4026_out0;
assign v$COUT_942_out0 = v$G1_4250_out0;
assign v$_10653_out0 = { v$_4551_out0,v$S_1250_out0 };
assign v$_10668_out0 = { v$_4566_out0,v$S_1474_out0 };
assign v$_10948_out0 = { v$_10653_out0,v$COUT_718_out0 };
assign v$_10963_out0 = { v$_10668_out0,v$COUT_942_out0 };
assign v$COUT_10918_out0 = v$_10948_out0;
assign v$COUT_10933_out0 = v$_10963_out0;
assign v$CIN_2359_out0 = v$COUT_10918_out0;
assign v$CIN_2374_out0 = v$COUT_10933_out0;
assign v$_472_out0 = v$CIN_2359_out0[8:8];
assign v$_487_out0 = v$CIN_2374_out0[8:8];
assign v$_1777_out0 = v$CIN_2359_out0[6:6];
assign v$_1792_out0 = v$CIN_2374_out0[6:6];
assign v$_2159_out0 = v$CIN_2359_out0[3:3];
assign v$_2174_out0 = v$CIN_2374_out0[3:3];
assign v$_2198_out0 = v$CIN_2359_out0[15:15];
assign v$_2212_out0 = v$CIN_2374_out0[15:15];
assign v$_2506_out0 = v$CIN_2359_out0[0:0];
assign v$_2521_out0 = v$CIN_2374_out0[0:0];
assign v$_3055_out0 = v$CIN_2359_out0[9:9];
assign v$_3070_out0 = v$CIN_2374_out0[9:9];
assign v$_3089_out0 = v$CIN_2359_out0[2:2];
assign v$_3104_out0 = v$CIN_2374_out0[2:2];
assign v$_3143_out0 = v$CIN_2359_out0[7:7];
assign v$_3158_out0 = v$CIN_2374_out0[7:7];
assign v$_3827_out0 = v$CIN_2359_out0[1:1];
assign v$_3842_out0 = v$CIN_2374_out0[1:1];
assign v$_3865_out0 = v$CIN_2359_out0[10:10];
assign v$_3880_out0 = v$CIN_2374_out0[10:10];
assign v$_6804_out0 = v$CIN_2359_out0[11:11];
assign v$_6819_out0 = v$CIN_2374_out0[11:11];
assign v$_7648_out0 = v$CIN_2359_out0[12:12];
assign v$_7663_out0 = v$CIN_2374_out0[12:12];
assign v$_8703_out0 = v$CIN_2359_out0[13:13];
assign v$_8718_out0 = v$CIN_2374_out0[13:13];
assign v$_8773_out0 = v$CIN_2359_out0[14:14];
assign v$_8788_out0 = v$CIN_2374_out0[14:14];
assign v$_10723_out0 = v$CIN_2359_out0[5:5];
assign v$_10738_out0 = v$CIN_2374_out0[5:5];
assign v$_13452_out0 = v$CIN_2359_out0[4:4];
assign v$_13467_out0 = v$CIN_2374_out0[4:4];
assign v$RM_3414_out0 = v$_7648_out0;
assign v$RM_3415_out0 = v$_8773_out0;
assign v$RM_3417_out0 = v$_10723_out0;
assign v$RM_3418_out0 = v$_13452_out0;
assign v$RM_3419_out0 = v$_8703_out0;
assign v$RM_3420_out0 = v$_3055_out0;
assign v$RM_3421_out0 = v$_3865_out0;
assign v$RM_3422_out0 = v$_3827_out0;
assign v$RM_3423_out0 = v$_2159_out0;
assign v$RM_3424_out0 = v$_1777_out0;
assign v$RM_3425_out0 = v$_3143_out0;
assign v$RM_3426_out0 = v$_6804_out0;
assign v$RM_3427_out0 = v$_472_out0;
assign v$RM_3428_out0 = v$_3089_out0;
assign v$RM_3638_out0 = v$_7663_out0;
assign v$RM_3639_out0 = v$_8788_out0;
assign v$RM_3641_out0 = v$_10738_out0;
assign v$RM_3642_out0 = v$_13467_out0;
assign v$RM_3643_out0 = v$_8718_out0;
assign v$RM_3644_out0 = v$_3070_out0;
assign v$RM_3645_out0 = v$_3880_out0;
assign v$RM_3646_out0 = v$_3842_out0;
assign v$RM_3647_out0 = v$_2174_out0;
assign v$RM_3648_out0 = v$_1792_out0;
assign v$RM_3649_out0 = v$_3158_out0;
assign v$RM_3650_out0 = v$_6819_out0;
assign v$RM_3651_out0 = v$_487_out0;
assign v$RM_3652_out0 = v$_3104_out0;
assign v$CIN_9869_out0 = v$_2198_out0;
assign v$CIN_10093_out0 = v$_2212_out0;
assign v$RM_11437_out0 = v$_2506_out0;
assign v$RM_11901_out0 = v$_2521_out0;
assign v$RD_5990_out0 = v$CIN_9869_out0;
assign v$RD_6454_out0 = v$CIN_10093_out0;
assign v$G1_7852_out0 = ((v$RD_5997_out0 && !v$RM_11437_out0) || (!v$RD_5997_out0) && v$RM_11437_out0);
assign v$G1_8316_out0 = ((v$RD_6461_out0 && !v$RM_11901_out0) || (!v$RD_6461_out0) && v$RM_11901_out0);
assign v$RM_11425_out0 = v$RM_3414_out0;
assign v$RM_11427_out0 = v$RM_3415_out0;
assign v$RM_11431_out0 = v$RM_3417_out0;
assign v$RM_11433_out0 = v$RM_3418_out0;
assign v$RM_11435_out0 = v$RM_3419_out0;
assign v$RM_11438_out0 = v$RM_3420_out0;
assign v$RM_11440_out0 = v$RM_3421_out0;
assign v$RM_11442_out0 = v$RM_3422_out0;
assign v$RM_11444_out0 = v$RM_3423_out0;
assign v$RM_11446_out0 = v$RM_3424_out0;
assign v$RM_11448_out0 = v$RM_3425_out0;
assign v$RM_11450_out0 = v$RM_3426_out0;
assign v$RM_11452_out0 = v$RM_3427_out0;
assign v$RM_11454_out0 = v$RM_3428_out0;
assign v$RM_11889_out0 = v$RM_3638_out0;
assign v$RM_11891_out0 = v$RM_3639_out0;
assign v$RM_11895_out0 = v$RM_3641_out0;
assign v$RM_11897_out0 = v$RM_3642_out0;
assign v$RM_11899_out0 = v$RM_3643_out0;
assign v$RM_11902_out0 = v$RM_3644_out0;
assign v$RM_11904_out0 = v$RM_3645_out0;
assign v$RM_11906_out0 = v$RM_3646_out0;
assign v$RM_11908_out0 = v$RM_3647_out0;
assign v$RM_11910_out0 = v$RM_3648_out0;
assign v$RM_11912_out0 = v$RM_3649_out0;
assign v$RM_11914_out0 = v$RM_3650_out0;
assign v$RM_11916_out0 = v$RM_3651_out0;
assign v$RM_11918_out0 = v$RM_3652_out0;
assign v$G2_12388_out0 = v$RD_5997_out0 && v$RM_11437_out0;
assign v$G2_12852_out0 = v$RD_6461_out0 && v$RM_11901_out0;
assign v$CARRY_4997_out0 = v$G2_12388_out0;
assign v$CARRY_5461_out0 = v$G2_12852_out0;
assign v$G1_7840_out0 = ((v$RD_5985_out0 && !v$RM_11425_out0) || (!v$RD_5985_out0) && v$RM_11425_out0);
assign v$G1_7842_out0 = ((v$RD_5987_out0 && !v$RM_11427_out0) || (!v$RD_5987_out0) && v$RM_11427_out0);
assign v$G1_7846_out0 = ((v$RD_5991_out0 && !v$RM_11431_out0) || (!v$RD_5991_out0) && v$RM_11431_out0);
assign v$G1_7848_out0 = ((v$RD_5993_out0 && !v$RM_11433_out0) || (!v$RD_5993_out0) && v$RM_11433_out0);
assign v$G1_7850_out0 = ((v$RD_5995_out0 && !v$RM_11435_out0) || (!v$RD_5995_out0) && v$RM_11435_out0);
assign v$G1_7853_out0 = ((v$RD_5998_out0 && !v$RM_11438_out0) || (!v$RD_5998_out0) && v$RM_11438_out0);
assign v$G1_7855_out0 = ((v$RD_6000_out0 && !v$RM_11440_out0) || (!v$RD_6000_out0) && v$RM_11440_out0);
assign v$G1_7857_out0 = ((v$RD_6002_out0 && !v$RM_11442_out0) || (!v$RD_6002_out0) && v$RM_11442_out0);
assign v$G1_7859_out0 = ((v$RD_6004_out0 && !v$RM_11444_out0) || (!v$RD_6004_out0) && v$RM_11444_out0);
assign v$G1_7861_out0 = ((v$RD_6006_out0 && !v$RM_11446_out0) || (!v$RD_6006_out0) && v$RM_11446_out0);
assign v$G1_7863_out0 = ((v$RD_6008_out0 && !v$RM_11448_out0) || (!v$RD_6008_out0) && v$RM_11448_out0);
assign v$G1_7865_out0 = ((v$RD_6010_out0 && !v$RM_11450_out0) || (!v$RD_6010_out0) && v$RM_11450_out0);
assign v$G1_7867_out0 = ((v$RD_6012_out0 && !v$RM_11452_out0) || (!v$RD_6012_out0) && v$RM_11452_out0);
assign v$G1_7869_out0 = ((v$RD_6014_out0 && !v$RM_11454_out0) || (!v$RD_6014_out0) && v$RM_11454_out0);
assign v$G1_8304_out0 = ((v$RD_6449_out0 && !v$RM_11889_out0) || (!v$RD_6449_out0) && v$RM_11889_out0);
assign v$G1_8306_out0 = ((v$RD_6451_out0 && !v$RM_11891_out0) || (!v$RD_6451_out0) && v$RM_11891_out0);
assign v$G1_8310_out0 = ((v$RD_6455_out0 && !v$RM_11895_out0) || (!v$RD_6455_out0) && v$RM_11895_out0);
assign v$G1_8312_out0 = ((v$RD_6457_out0 && !v$RM_11897_out0) || (!v$RD_6457_out0) && v$RM_11897_out0);
assign v$G1_8314_out0 = ((v$RD_6459_out0 && !v$RM_11899_out0) || (!v$RD_6459_out0) && v$RM_11899_out0);
assign v$G1_8317_out0 = ((v$RD_6462_out0 && !v$RM_11902_out0) || (!v$RD_6462_out0) && v$RM_11902_out0);
assign v$G1_8319_out0 = ((v$RD_6464_out0 && !v$RM_11904_out0) || (!v$RD_6464_out0) && v$RM_11904_out0);
assign v$G1_8321_out0 = ((v$RD_6466_out0 && !v$RM_11906_out0) || (!v$RD_6466_out0) && v$RM_11906_out0);
assign v$G1_8323_out0 = ((v$RD_6468_out0 && !v$RM_11908_out0) || (!v$RD_6468_out0) && v$RM_11908_out0);
assign v$G1_8325_out0 = ((v$RD_6470_out0 && !v$RM_11910_out0) || (!v$RD_6470_out0) && v$RM_11910_out0);
assign v$G1_8327_out0 = ((v$RD_6472_out0 && !v$RM_11912_out0) || (!v$RD_6472_out0) && v$RM_11912_out0);
assign v$G1_8329_out0 = ((v$RD_6474_out0 && !v$RM_11914_out0) || (!v$RD_6474_out0) && v$RM_11914_out0);
assign v$G1_8331_out0 = ((v$RD_6476_out0 && !v$RM_11916_out0) || (!v$RD_6476_out0) && v$RM_11916_out0);
assign v$G1_8333_out0 = ((v$RD_6478_out0 && !v$RM_11918_out0) || (!v$RD_6478_out0) && v$RM_11918_out0);
assign v$S_8998_out0 = v$G1_7852_out0;
assign v$S_9462_out0 = v$G1_8316_out0;
assign v$G2_12376_out0 = v$RD_5985_out0 && v$RM_11425_out0;
assign v$G2_12378_out0 = v$RD_5987_out0 && v$RM_11427_out0;
assign v$G2_12382_out0 = v$RD_5991_out0 && v$RM_11431_out0;
assign v$G2_12384_out0 = v$RD_5993_out0 && v$RM_11433_out0;
assign v$G2_12386_out0 = v$RD_5995_out0 && v$RM_11435_out0;
assign v$G2_12389_out0 = v$RD_5998_out0 && v$RM_11438_out0;
assign v$G2_12391_out0 = v$RD_6000_out0 && v$RM_11440_out0;
assign v$G2_12393_out0 = v$RD_6002_out0 && v$RM_11442_out0;
assign v$G2_12395_out0 = v$RD_6004_out0 && v$RM_11444_out0;
assign v$G2_12397_out0 = v$RD_6006_out0 && v$RM_11446_out0;
assign v$G2_12399_out0 = v$RD_6008_out0 && v$RM_11448_out0;
assign v$G2_12401_out0 = v$RD_6010_out0 && v$RM_11450_out0;
assign v$G2_12403_out0 = v$RD_6012_out0 && v$RM_11452_out0;
assign v$G2_12405_out0 = v$RD_6014_out0 && v$RM_11454_out0;
assign v$G2_12840_out0 = v$RD_6449_out0 && v$RM_11889_out0;
assign v$G2_12842_out0 = v$RD_6451_out0 && v$RM_11891_out0;
assign v$G2_12846_out0 = v$RD_6455_out0 && v$RM_11895_out0;
assign v$G2_12848_out0 = v$RD_6457_out0 && v$RM_11897_out0;
assign v$G2_12850_out0 = v$RD_6459_out0 && v$RM_11899_out0;
assign v$G2_12853_out0 = v$RD_6462_out0 && v$RM_11902_out0;
assign v$G2_12855_out0 = v$RD_6464_out0 && v$RM_11904_out0;
assign v$G2_12857_out0 = v$RD_6466_out0 && v$RM_11906_out0;
assign v$G2_12859_out0 = v$RD_6468_out0 && v$RM_11908_out0;
assign v$G2_12861_out0 = v$RD_6470_out0 && v$RM_11910_out0;
assign v$G2_12863_out0 = v$RD_6472_out0 && v$RM_11912_out0;
assign v$G2_12865_out0 = v$RD_6474_out0 && v$RM_11914_out0;
assign v$G2_12867_out0 = v$RD_6476_out0 && v$RM_11916_out0;
assign v$G2_12869_out0 = v$RD_6478_out0 && v$RM_11918_out0;
assign v$S_4669_out0 = v$S_8998_out0;
assign v$S_4684_out0 = v$S_9462_out0;
assign v$CARRY_4985_out0 = v$G2_12376_out0;
assign v$CARRY_4987_out0 = v$G2_12378_out0;
assign v$CARRY_4991_out0 = v$G2_12382_out0;
assign v$CARRY_4993_out0 = v$G2_12384_out0;
assign v$CARRY_4995_out0 = v$G2_12386_out0;
assign v$CARRY_4998_out0 = v$G2_12389_out0;
assign v$CARRY_5000_out0 = v$G2_12391_out0;
assign v$CARRY_5002_out0 = v$G2_12393_out0;
assign v$CARRY_5004_out0 = v$G2_12395_out0;
assign v$CARRY_5006_out0 = v$G2_12397_out0;
assign v$CARRY_5008_out0 = v$G2_12399_out0;
assign v$CARRY_5010_out0 = v$G2_12401_out0;
assign v$CARRY_5012_out0 = v$G2_12403_out0;
assign v$CARRY_5014_out0 = v$G2_12405_out0;
assign v$CARRY_5449_out0 = v$G2_12840_out0;
assign v$CARRY_5451_out0 = v$G2_12842_out0;
assign v$CARRY_5455_out0 = v$G2_12846_out0;
assign v$CARRY_5457_out0 = v$G2_12848_out0;
assign v$CARRY_5459_out0 = v$G2_12850_out0;
assign v$CARRY_5462_out0 = v$G2_12853_out0;
assign v$CARRY_5464_out0 = v$G2_12855_out0;
assign v$CARRY_5466_out0 = v$G2_12857_out0;
assign v$CARRY_5468_out0 = v$G2_12859_out0;
assign v$CARRY_5470_out0 = v$G2_12861_out0;
assign v$CARRY_5472_out0 = v$G2_12863_out0;
assign v$CARRY_5474_out0 = v$G2_12865_out0;
assign v$CARRY_5476_out0 = v$G2_12867_out0;
assign v$CARRY_5478_out0 = v$G2_12869_out0;
assign v$S_8986_out0 = v$G1_7840_out0;
assign v$S_8988_out0 = v$G1_7842_out0;
assign v$S_8992_out0 = v$G1_7846_out0;
assign v$S_8994_out0 = v$G1_7848_out0;
assign v$S_8996_out0 = v$G1_7850_out0;
assign v$S_8999_out0 = v$G1_7853_out0;
assign v$S_9001_out0 = v$G1_7855_out0;
assign v$S_9003_out0 = v$G1_7857_out0;
assign v$S_9005_out0 = v$G1_7859_out0;
assign v$S_9007_out0 = v$G1_7861_out0;
assign v$S_9009_out0 = v$G1_7863_out0;
assign v$S_9011_out0 = v$G1_7865_out0;
assign v$S_9013_out0 = v$G1_7867_out0;
assign v$S_9015_out0 = v$G1_7869_out0;
assign v$S_9450_out0 = v$G1_8304_out0;
assign v$S_9452_out0 = v$G1_8306_out0;
assign v$S_9456_out0 = v$G1_8310_out0;
assign v$S_9458_out0 = v$G1_8312_out0;
assign v$S_9460_out0 = v$G1_8314_out0;
assign v$S_9463_out0 = v$G1_8317_out0;
assign v$S_9465_out0 = v$G1_8319_out0;
assign v$S_9467_out0 = v$G1_8321_out0;
assign v$S_9469_out0 = v$G1_8323_out0;
assign v$S_9471_out0 = v$G1_8325_out0;
assign v$S_9473_out0 = v$G1_8327_out0;
assign v$S_9475_out0 = v$G1_8329_out0;
assign v$S_9477_out0 = v$G1_8331_out0;
assign v$S_9479_out0 = v$G1_8333_out0;
assign v$CIN_9875_out0 = v$CARRY_4997_out0;
assign v$CIN_10099_out0 = v$CARRY_5461_out0;
assign v$_4529_out0 = { v$_1716_out0,v$S_4669_out0 };
assign v$_4530_out0 = { v$_1717_out0,v$S_4684_out0 };
assign v$RD_6003_out0 = v$CIN_9875_out0;
assign v$RD_6467_out0 = v$CIN_10099_out0;
assign v$RM_11426_out0 = v$S_8986_out0;
assign v$RM_11428_out0 = v$S_8988_out0;
assign v$RM_11432_out0 = v$S_8992_out0;
assign v$RM_11434_out0 = v$S_8994_out0;
assign v$RM_11436_out0 = v$S_8996_out0;
assign v$RM_11439_out0 = v$S_8999_out0;
assign v$RM_11441_out0 = v$S_9001_out0;
assign v$RM_11443_out0 = v$S_9003_out0;
assign v$RM_11445_out0 = v$S_9005_out0;
assign v$RM_11447_out0 = v$S_9007_out0;
assign v$RM_11449_out0 = v$S_9009_out0;
assign v$RM_11451_out0 = v$S_9011_out0;
assign v$RM_11453_out0 = v$S_9013_out0;
assign v$RM_11455_out0 = v$S_9015_out0;
assign v$RM_11890_out0 = v$S_9450_out0;
assign v$RM_11892_out0 = v$S_9452_out0;
assign v$RM_11896_out0 = v$S_9456_out0;
assign v$RM_11898_out0 = v$S_9458_out0;
assign v$RM_11900_out0 = v$S_9460_out0;
assign v$RM_11903_out0 = v$S_9463_out0;
assign v$RM_11905_out0 = v$S_9465_out0;
assign v$RM_11907_out0 = v$S_9467_out0;
assign v$RM_11909_out0 = v$S_9469_out0;
assign v$RM_11911_out0 = v$S_9471_out0;
assign v$RM_11913_out0 = v$S_9473_out0;
assign v$RM_11915_out0 = v$S_9475_out0;
assign v$RM_11917_out0 = v$S_9477_out0;
assign v$RM_11919_out0 = v$S_9479_out0;
assign v$G1_7858_out0 = ((v$RD_6003_out0 && !v$RM_11443_out0) || (!v$RD_6003_out0) && v$RM_11443_out0);
assign v$G1_8322_out0 = ((v$RD_6467_out0 && !v$RM_11907_out0) || (!v$RD_6467_out0) && v$RM_11907_out0);
assign v$G2_12394_out0 = v$RD_6003_out0 && v$RM_11443_out0;
assign v$G2_12858_out0 = v$RD_6467_out0 && v$RM_11907_out0;
assign v$CARRY_5003_out0 = v$G2_12394_out0;
assign v$CARRY_5467_out0 = v$G2_12858_out0;
assign v$S_9004_out0 = v$G1_7858_out0;
assign v$S_9468_out0 = v$G1_8322_out0;
assign v$S_1286_out0 = v$S_9004_out0;
assign v$S_1510_out0 = v$S_9468_out0;
assign v$G1_4062_out0 = v$CARRY_5003_out0 || v$CARRY_5002_out0;
assign v$G1_4286_out0 = v$CARRY_5467_out0 || v$CARRY_5466_out0;
assign v$COUT_754_out0 = v$G1_4062_out0;
assign v$COUT_978_out0 = v$G1_4286_out0;
assign v$CIN_9881_out0 = v$COUT_754_out0;
assign v$CIN_10105_out0 = v$COUT_978_out0;
assign v$RD_6015_out0 = v$CIN_9881_out0;
assign v$RD_6479_out0 = v$CIN_10105_out0;
assign v$G1_7870_out0 = ((v$RD_6015_out0 && !v$RM_11455_out0) || (!v$RD_6015_out0) && v$RM_11455_out0);
assign v$G1_8334_out0 = ((v$RD_6479_out0 && !v$RM_11919_out0) || (!v$RD_6479_out0) && v$RM_11919_out0);
assign v$G2_12406_out0 = v$RD_6015_out0 && v$RM_11455_out0;
assign v$G2_12870_out0 = v$RD_6479_out0 && v$RM_11919_out0;
assign v$CARRY_5015_out0 = v$G2_12406_out0;
assign v$CARRY_5479_out0 = v$G2_12870_out0;
assign v$S_9016_out0 = v$G1_7870_out0;
assign v$S_9480_out0 = v$G1_8334_out0;
assign v$S_1292_out0 = v$S_9016_out0;
assign v$S_1516_out0 = v$S_9480_out0;
assign v$G1_4068_out0 = v$CARRY_5015_out0 || v$CARRY_5014_out0;
assign v$G1_4292_out0 = v$CARRY_5479_out0 || v$CARRY_5478_out0;
assign v$COUT_760_out0 = v$G1_4068_out0;
assign v$COUT_984_out0 = v$G1_4292_out0;
assign v$_4786_out0 = { v$S_1286_out0,v$S_1292_out0 };
assign v$_4801_out0 = { v$S_1510_out0,v$S_1516_out0 };
assign v$CIN_9876_out0 = v$COUT_760_out0;
assign v$CIN_10100_out0 = v$COUT_984_out0;
assign v$RD_6005_out0 = v$CIN_9876_out0;
assign v$RD_6469_out0 = v$CIN_10100_out0;
assign v$G1_7860_out0 = ((v$RD_6005_out0 && !v$RM_11445_out0) || (!v$RD_6005_out0) && v$RM_11445_out0);
assign v$G1_8324_out0 = ((v$RD_6469_out0 && !v$RM_11909_out0) || (!v$RD_6469_out0) && v$RM_11909_out0);
assign v$G2_12396_out0 = v$RD_6005_out0 && v$RM_11445_out0;
assign v$G2_12860_out0 = v$RD_6469_out0 && v$RM_11909_out0;
assign v$CARRY_5005_out0 = v$G2_12396_out0;
assign v$CARRY_5469_out0 = v$G2_12860_out0;
assign v$S_9006_out0 = v$G1_7860_out0;
assign v$S_9470_out0 = v$G1_8324_out0;
assign v$S_1287_out0 = v$S_9006_out0;
assign v$S_1511_out0 = v$S_9470_out0;
assign v$G1_4063_out0 = v$CARRY_5005_out0 || v$CARRY_5004_out0;
assign v$G1_4287_out0 = v$CARRY_5469_out0 || v$CARRY_5468_out0;
assign v$COUT_755_out0 = v$G1_4063_out0;
assign v$COUT_979_out0 = v$G1_4287_out0;
assign v$_2556_out0 = { v$_4786_out0,v$S_1287_out0 };
assign v$_2571_out0 = { v$_4801_out0,v$S_1511_out0 };
assign v$CIN_9871_out0 = v$COUT_755_out0;
assign v$CIN_10095_out0 = v$COUT_979_out0;
assign v$RD_5994_out0 = v$CIN_9871_out0;
assign v$RD_6458_out0 = v$CIN_10095_out0;
assign v$G1_7849_out0 = ((v$RD_5994_out0 && !v$RM_11434_out0) || (!v$RD_5994_out0) && v$RM_11434_out0);
assign v$G1_8313_out0 = ((v$RD_6458_out0 && !v$RM_11898_out0) || (!v$RD_6458_out0) && v$RM_11898_out0);
assign v$G2_12385_out0 = v$RD_5994_out0 && v$RM_11434_out0;
assign v$G2_12849_out0 = v$RD_6458_out0 && v$RM_11898_out0;
assign v$CARRY_4994_out0 = v$G2_12385_out0;
assign v$CARRY_5458_out0 = v$G2_12849_out0;
assign v$S_8995_out0 = v$G1_7849_out0;
assign v$S_9459_out0 = v$G1_8313_out0;
assign v$S_1282_out0 = v$S_8995_out0;
assign v$S_1506_out0 = v$S_9459_out0;
assign v$G1_4058_out0 = v$CARRY_4994_out0 || v$CARRY_4993_out0;
assign v$G1_4282_out0 = v$CARRY_5458_out0 || v$CARRY_5457_out0;
assign v$COUT_750_out0 = v$G1_4058_out0;
assign v$COUT_974_out0 = v$G1_4282_out0;
assign v$_7036_out0 = { v$_2556_out0,v$S_1282_out0 };
assign v$_7051_out0 = { v$_2571_out0,v$S_1506_out0 };
assign v$CIN_9870_out0 = v$COUT_750_out0;
assign v$CIN_10094_out0 = v$COUT_974_out0;
assign v$RD_5992_out0 = v$CIN_9870_out0;
assign v$RD_6456_out0 = v$CIN_10094_out0;
assign v$G1_7847_out0 = ((v$RD_5992_out0 && !v$RM_11432_out0) || (!v$RD_5992_out0) && v$RM_11432_out0);
assign v$G1_8311_out0 = ((v$RD_6456_out0 && !v$RM_11896_out0) || (!v$RD_6456_out0) && v$RM_11896_out0);
assign v$G2_12383_out0 = v$RD_5992_out0 && v$RM_11432_out0;
assign v$G2_12847_out0 = v$RD_6456_out0 && v$RM_11896_out0;
assign v$CARRY_4992_out0 = v$G2_12383_out0;
assign v$CARRY_5456_out0 = v$G2_12847_out0;
assign v$S_8993_out0 = v$G1_7847_out0;
assign v$S_9457_out0 = v$G1_8311_out0;
assign v$S_1281_out0 = v$S_8993_out0;
assign v$S_1505_out0 = v$S_9457_out0;
assign v$G1_4057_out0 = v$CARRY_4992_out0 || v$CARRY_4991_out0;
assign v$G1_4281_out0 = v$CARRY_5456_out0 || v$CARRY_5455_out0;
assign v$COUT_749_out0 = v$G1_4057_out0;
assign v$COUT_973_out0 = v$G1_4281_out0;
assign v$_13522_out0 = { v$_7036_out0,v$S_1281_out0 };
assign v$_13537_out0 = { v$_7051_out0,v$S_1505_out0 };
assign v$CIN_9877_out0 = v$COUT_749_out0;
assign v$CIN_10101_out0 = v$COUT_973_out0;
assign v$RD_6007_out0 = v$CIN_9877_out0;
assign v$RD_6471_out0 = v$CIN_10101_out0;
assign v$G1_7862_out0 = ((v$RD_6007_out0 && !v$RM_11447_out0) || (!v$RD_6007_out0) && v$RM_11447_out0);
assign v$G1_8326_out0 = ((v$RD_6471_out0 && !v$RM_11911_out0) || (!v$RD_6471_out0) && v$RM_11911_out0);
assign v$G2_12398_out0 = v$RD_6007_out0 && v$RM_11447_out0;
assign v$G2_12862_out0 = v$RD_6471_out0 && v$RM_11911_out0;
assign v$CARRY_5007_out0 = v$G2_12398_out0;
assign v$CARRY_5471_out0 = v$G2_12862_out0;
assign v$S_9008_out0 = v$G1_7862_out0;
assign v$S_9472_out0 = v$G1_8326_out0;
assign v$S_1288_out0 = v$S_9008_out0;
assign v$S_1512_out0 = v$S_9472_out0;
assign v$G1_4064_out0 = v$CARRY_5007_out0 || v$CARRY_5006_out0;
assign v$G1_4288_out0 = v$CARRY_5471_out0 || v$CARRY_5470_out0;
assign v$COUT_756_out0 = v$G1_4064_out0;
assign v$COUT_980_out0 = v$G1_4288_out0;
assign v$_3315_out0 = { v$_13522_out0,v$S_1288_out0 };
assign v$_3330_out0 = { v$_13537_out0,v$S_1512_out0 };
assign v$CIN_9878_out0 = v$COUT_756_out0;
assign v$CIN_10102_out0 = v$COUT_980_out0;
assign v$RD_6009_out0 = v$CIN_9878_out0;
assign v$RD_6473_out0 = v$CIN_10102_out0;
assign v$G1_7864_out0 = ((v$RD_6009_out0 && !v$RM_11449_out0) || (!v$RD_6009_out0) && v$RM_11449_out0);
assign v$G1_8328_out0 = ((v$RD_6473_out0 && !v$RM_11913_out0) || (!v$RD_6473_out0) && v$RM_11913_out0);
assign v$G2_12400_out0 = v$RD_6009_out0 && v$RM_11449_out0;
assign v$G2_12864_out0 = v$RD_6473_out0 && v$RM_11913_out0;
assign v$CARRY_5009_out0 = v$G2_12400_out0;
assign v$CARRY_5473_out0 = v$G2_12864_out0;
assign v$S_9010_out0 = v$G1_7864_out0;
assign v$S_9474_out0 = v$G1_8328_out0;
assign v$S_1289_out0 = v$S_9010_out0;
assign v$S_1513_out0 = v$S_9474_out0;
assign v$G1_4065_out0 = v$CARRY_5009_out0 || v$CARRY_5008_out0;
assign v$G1_4289_out0 = v$CARRY_5473_out0 || v$CARRY_5472_out0;
assign v$COUT_757_out0 = v$G1_4065_out0;
assign v$COUT_981_out0 = v$G1_4289_out0;
assign v$_7151_out0 = { v$_3315_out0,v$S_1289_out0 };
assign v$_7166_out0 = { v$_3330_out0,v$S_1513_out0 };
assign v$CIN_9880_out0 = v$COUT_757_out0;
assign v$CIN_10104_out0 = v$COUT_981_out0;
assign v$RD_6013_out0 = v$CIN_9880_out0;
assign v$RD_6477_out0 = v$CIN_10104_out0;
assign v$G1_7868_out0 = ((v$RD_6013_out0 && !v$RM_11453_out0) || (!v$RD_6013_out0) && v$RM_11453_out0);
assign v$G1_8332_out0 = ((v$RD_6477_out0 && !v$RM_11917_out0) || (!v$RD_6477_out0) && v$RM_11917_out0);
assign v$G2_12404_out0 = v$RD_6013_out0 && v$RM_11453_out0;
assign v$G2_12868_out0 = v$RD_6477_out0 && v$RM_11917_out0;
assign v$CARRY_5013_out0 = v$G2_12404_out0;
assign v$CARRY_5477_out0 = v$G2_12868_out0;
assign v$S_9014_out0 = v$G1_7868_out0;
assign v$S_9478_out0 = v$G1_8332_out0;
assign v$S_1291_out0 = v$S_9014_out0;
assign v$S_1515_out0 = v$S_9478_out0;
assign v$G1_4067_out0 = v$CARRY_5013_out0 || v$CARRY_5012_out0;
assign v$G1_4291_out0 = v$CARRY_5477_out0 || v$CARRY_5476_out0;
assign v$COUT_759_out0 = v$G1_4067_out0;
assign v$COUT_983_out0 = v$G1_4291_out0;
assign v$_4753_out0 = { v$_7151_out0,v$S_1291_out0 };
assign v$_4768_out0 = { v$_7166_out0,v$S_1515_out0 };
assign v$CIN_9873_out0 = v$COUT_759_out0;
assign v$CIN_10097_out0 = v$COUT_983_out0;
assign v$RD_5999_out0 = v$CIN_9873_out0;
assign v$RD_6463_out0 = v$CIN_10097_out0;
assign v$G1_7854_out0 = ((v$RD_5999_out0 && !v$RM_11439_out0) || (!v$RD_5999_out0) && v$RM_11439_out0);
assign v$G1_8318_out0 = ((v$RD_6463_out0 && !v$RM_11903_out0) || (!v$RD_6463_out0) && v$RM_11903_out0);
assign v$G2_12390_out0 = v$RD_5999_out0 && v$RM_11439_out0;
assign v$G2_12854_out0 = v$RD_6463_out0 && v$RM_11903_out0;
assign v$CARRY_4999_out0 = v$G2_12390_out0;
assign v$CARRY_5463_out0 = v$G2_12854_out0;
assign v$S_9000_out0 = v$G1_7854_out0;
assign v$S_9464_out0 = v$G1_8318_out0;
assign v$S_1284_out0 = v$S_9000_out0;
assign v$S_1508_out0 = v$S_9464_out0;
assign v$G1_4060_out0 = v$CARRY_4999_out0 || v$CARRY_4998_out0;
assign v$G1_4284_out0 = v$CARRY_5463_out0 || v$CARRY_5462_out0;
assign v$COUT_752_out0 = v$G1_4060_out0;
assign v$COUT_976_out0 = v$G1_4284_out0;
assign v$_6930_out0 = { v$_4753_out0,v$S_1284_out0 };
assign v$_6945_out0 = { v$_4768_out0,v$S_1508_out0 };
assign v$CIN_9874_out0 = v$COUT_752_out0;
assign v$CIN_10098_out0 = v$COUT_976_out0;
assign v$RD_6001_out0 = v$CIN_9874_out0;
assign v$RD_6465_out0 = v$CIN_10098_out0;
assign v$G1_7856_out0 = ((v$RD_6001_out0 && !v$RM_11441_out0) || (!v$RD_6001_out0) && v$RM_11441_out0);
assign v$G1_8320_out0 = ((v$RD_6465_out0 && !v$RM_11905_out0) || (!v$RD_6465_out0) && v$RM_11905_out0);
assign v$G2_12392_out0 = v$RD_6001_out0 && v$RM_11441_out0;
assign v$G2_12856_out0 = v$RD_6465_out0 && v$RM_11905_out0;
assign v$CARRY_5001_out0 = v$G2_12392_out0;
assign v$CARRY_5465_out0 = v$G2_12856_out0;
assign v$S_9002_out0 = v$G1_7856_out0;
assign v$S_9466_out0 = v$G1_8320_out0;
assign v$S_1285_out0 = v$S_9002_out0;
assign v$S_1509_out0 = v$S_9466_out0;
assign v$G1_4061_out0 = v$CARRY_5001_out0 || v$CARRY_5000_out0;
assign v$G1_4285_out0 = v$CARRY_5465_out0 || v$CARRY_5464_out0;
assign v$COUT_753_out0 = v$G1_4061_out0;
assign v$COUT_977_out0 = v$G1_4285_out0;
assign v$_5806_out0 = { v$_6930_out0,v$S_1285_out0 };
assign v$_5821_out0 = { v$_6945_out0,v$S_1509_out0 };
assign v$CIN_9879_out0 = v$COUT_753_out0;
assign v$CIN_10103_out0 = v$COUT_977_out0;
assign v$RD_6011_out0 = v$CIN_9879_out0;
assign v$RD_6475_out0 = v$CIN_10103_out0;
assign v$G1_7866_out0 = ((v$RD_6011_out0 && !v$RM_11451_out0) || (!v$RD_6011_out0) && v$RM_11451_out0);
assign v$G1_8330_out0 = ((v$RD_6475_out0 && !v$RM_11915_out0) || (!v$RD_6475_out0) && v$RM_11915_out0);
assign v$G2_12402_out0 = v$RD_6011_out0 && v$RM_11451_out0;
assign v$G2_12866_out0 = v$RD_6475_out0 && v$RM_11915_out0;
assign v$CARRY_5011_out0 = v$G2_12402_out0;
assign v$CARRY_5475_out0 = v$G2_12866_out0;
assign v$S_9012_out0 = v$G1_7866_out0;
assign v$S_9476_out0 = v$G1_8330_out0;
assign v$S_1290_out0 = v$S_9012_out0;
assign v$S_1514_out0 = v$S_9476_out0;
assign v$G1_4066_out0 = v$CARRY_5011_out0 || v$CARRY_5010_out0;
assign v$G1_4290_out0 = v$CARRY_5475_out0 || v$CARRY_5474_out0;
assign v$COUT_758_out0 = v$G1_4066_out0;
assign v$COUT_982_out0 = v$G1_4290_out0;
assign v$_2030_out0 = { v$_5806_out0,v$S_1290_out0 };
assign v$_2045_out0 = { v$_5821_out0,v$S_1514_out0 };
assign v$CIN_9867_out0 = v$COUT_758_out0;
assign v$CIN_10091_out0 = v$COUT_982_out0;
assign v$RD_5986_out0 = v$CIN_9867_out0;
assign v$RD_6450_out0 = v$CIN_10091_out0;
assign v$G1_7841_out0 = ((v$RD_5986_out0 && !v$RM_11426_out0) || (!v$RD_5986_out0) && v$RM_11426_out0);
assign v$G1_8305_out0 = ((v$RD_6450_out0 && !v$RM_11890_out0) || (!v$RD_6450_out0) && v$RM_11890_out0);
assign v$G2_12377_out0 = v$RD_5986_out0 && v$RM_11426_out0;
assign v$G2_12841_out0 = v$RD_6450_out0 && v$RM_11890_out0;
assign v$CARRY_4986_out0 = v$G2_12377_out0;
assign v$CARRY_5450_out0 = v$G2_12841_out0;
assign v$S_8987_out0 = v$G1_7841_out0;
assign v$S_9451_out0 = v$G1_8305_out0;
assign v$S_1278_out0 = v$S_8987_out0;
assign v$S_1502_out0 = v$S_9451_out0;
assign v$G1_4054_out0 = v$CARRY_4986_out0 || v$CARRY_4985_out0;
assign v$G1_4278_out0 = v$CARRY_5450_out0 || v$CARRY_5449_out0;
assign v$COUT_746_out0 = v$G1_4054_out0;
assign v$COUT_970_out0 = v$G1_4278_out0;
assign v$_2797_out0 = { v$_2030_out0,v$S_1278_out0 };
assign v$_2812_out0 = { v$_2045_out0,v$S_1502_out0 };
assign v$CIN_9872_out0 = v$COUT_746_out0;
assign v$CIN_10096_out0 = v$COUT_970_out0;
assign v$RD_5996_out0 = v$CIN_9872_out0;
assign v$RD_6460_out0 = v$CIN_10096_out0;
assign v$G1_7851_out0 = ((v$RD_5996_out0 && !v$RM_11436_out0) || (!v$RD_5996_out0) && v$RM_11436_out0);
assign v$G1_8315_out0 = ((v$RD_6460_out0 && !v$RM_11900_out0) || (!v$RD_6460_out0) && v$RM_11900_out0);
assign v$G2_12387_out0 = v$RD_5996_out0 && v$RM_11436_out0;
assign v$G2_12851_out0 = v$RD_6460_out0 && v$RM_11900_out0;
assign v$CARRY_4996_out0 = v$G2_12387_out0;
assign v$CARRY_5460_out0 = v$G2_12851_out0;
assign v$S_8997_out0 = v$G1_7851_out0;
assign v$S_9461_out0 = v$G1_8315_out0;
assign v$S_1283_out0 = v$S_8997_out0;
assign v$S_1507_out0 = v$S_9461_out0;
assign v$G1_4059_out0 = v$CARRY_4996_out0 || v$CARRY_4995_out0;
assign v$G1_4283_out0 = v$CARRY_5460_out0 || v$CARRY_5459_out0;
assign v$COUT_751_out0 = v$G1_4059_out0;
assign v$COUT_975_out0 = v$G1_4283_out0;
assign v$_1829_out0 = { v$_2797_out0,v$S_1283_out0 };
assign v$_1844_out0 = { v$_2812_out0,v$S_1507_out0 };
assign v$CIN_9868_out0 = v$COUT_751_out0;
assign v$CIN_10092_out0 = v$COUT_975_out0;
assign v$RD_5988_out0 = v$CIN_9868_out0;
assign v$RD_6452_out0 = v$CIN_10092_out0;
assign v$G1_7843_out0 = ((v$RD_5988_out0 && !v$RM_11428_out0) || (!v$RD_5988_out0) && v$RM_11428_out0);
assign v$G1_8307_out0 = ((v$RD_6452_out0 && !v$RM_11892_out0) || (!v$RD_6452_out0) && v$RM_11892_out0);
assign v$G2_12379_out0 = v$RD_5988_out0 && v$RM_11428_out0;
assign v$G2_12843_out0 = v$RD_6452_out0 && v$RM_11892_out0;
assign v$CARRY_4988_out0 = v$G2_12379_out0;
assign v$CARRY_5452_out0 = v$G2_12843_out0;
assign v$S_8989_out0 = v$G1_7843_out0;
assign v$S_9453_out0 = v$G1_8307_out0;
assign v$S_1279_out0 = v$S_8989_out0;
assign v$S_1503_out0 = v$S_9453_out0;
assign v$G1_4055_out0 = v$CARRY_4988_out0 || v$CARRY_4987_out0;
assign v$G1_4279_out0 = v$CARRY_5452_out0 || v$CARRY_5451_out0;
assign v$COUT_747_out0 = v$G1_4055_out0;
assign v$COUT_971_out0 = v$G1_4279_out0;
assign v$_4553_out0 = { v$_1829_out0,v$S_1279_out0 };
assign v$_4568_out0 = { v$_1844_out0,v$S_1503_out0 };
assign v$RM_3416_out0 = v$COUT_747_out0;
assign v$RM_3640_out0 = v$COUT_971_out0;
assign v$RM_11429_out0 = v$RM_3416_out0;
assign v$RM_11893_out0 = v$RM_3640_out0;
assign v$G1_7844_out0 = ((v$RD_5989_out0 && !v$RM_11429_out0) || (!v$RD_5989_out0) && v$RM_11429_out0);
assign v$G1_8308_out0 = ((v$RD_6453_out0 && !v$RM_11893_out0) || (!v$RD_6453_out0) && v$RM_11893_out0);
assign v$G2_12380_out0 = v$RD_5989_out0 && v$RM_11429_out0;
assign v$G2_12844_out0 = v$RD_6453_out0 && v$RM_11893_out0;
assign v$CARRY_4989_out0 = v$G2_12380_out0;
assign v$CARRY_5453_out0 = v$G2_12844_out0;
assign v$S_8990_out0 = v$G1_7844_out0;
assign v$S_9454_out0 = v$G1_8308_out0;
assign v$RM_11430_out0 = v$S_8990_out0;
assign v$RM_11894_out0 = v$S_9454_out0;
assign v$G1_7845_out0 = ((v$RD_5990_out0 && !v$RM_11430_out0) || (!v$RD_5990_out0) && v$RM_11430_out0);
assign v$G1_8309_out0 = ((v$RD_6454_out0 && !v$RM_11894_out0) || (!v$RD_6454_out0) && v$RM_11894_out0);
assign v$G2_12381_out0 = v$RD_5990_out0 && v$RM_11430_out0;
assign v$G2_12845_out0 = v$RD_6454_out0 && v$RM_11894_out0;
assign v$CARRY_4990_out0 = v$G2_12381_out0;
assign v$CARRY_5454_out0 = v$G2_12845_out0;
assign v$S_8991_out0 = v$G1_7845_out0;
assign v$S_9455_out0 = v$G1_8309_out0;
assign v$S_1280_out0 = v$S_8991_out0;
assign v$S_1504_out0 = v$S_9455_out0;
assign v$G1_4056_out0 = v$CARRY_4990_out0 || v$CARRY_4989_out0;
assign v$G1_4280_out0 = v$CARRY_5454_out0 || v$CARRY_5453_out0;
assign v$COUT_748_out0 = v$G1_4056_out0;
assign v$COUT_972_out0 = v$G1_4280_out0;
assign v$_10655_out0 = { v$_4553_out0,v$S_1280_out0 };
assign v$_10670_out0 = { v$_4568_out0,v$S_1504_out0 };
assign v$_10950_out0 = { v$_10655_out0,v$COUT_748_out0 };
assign v$_10965_out0 = { v$_10670_out0,v$COUT_972_out0 };
assign v$COUT_10920_out0 = v$_10950_out0;
assign v$COUT_10935_out0 = v$_10965_out0;
assign v$CIN_2355_out0 = v$COUT_10920_out0;
assign v$CIN_2370_out0 = v$COUT_10935_out0;
assign v$_468_out0 = v$CIN_2355_out0[8:8];
assign v$_483_out0 = v$CIN_2370_out0[8:8];
assign v$_1773_out0 = v$CIN_2355_out0[6:6];
assign v$_1788_out0 = v$CIN_2370_out0[6:6];
assign v$_2155_out0 = v$CIN_2355_out0[3:3];
assign v$_2170_out0 = v$CIN_2370_out0[3:3];
assign v$_2195_out0 = v$CIN_2355_out0[15:15];
assign v$_2209_out0 = v$CIN_2370_out0[15:15];
assign v$_2502_out0 = v$CIN_2355_out0[0:0];
assign v$_2517_out0 = v$CIN_2370_out0[0:0];
assign v$_3051_out0 = v$CIN_2355_out0[9:9];
assign v$_3066_out0 = v$CIN_2370_out0[9:9];
assign v$_3085_out0 = v$CIN_2355_out0[2:2];
assign v$_3100_out0 = v$CIN_2370_out0[2:2];
assign v$_3139_out0 = v$CIN_2355_out0[7:7];
assign v$_3154_out0 = v$CIN_2370_out0[7:7];
assign v$_3823_out0 = v$CIN_2355_out0[1:1];
assign v$_3838_out0 = v$CIN_2370_out0[1:1];
assign v$_3861_out0 = v$CIN_2355_out0[10:10];
assign v$_3876_out0 = v$CIN_2370_out0[10:10];
assign v$_6800_out0 = v$CIN_2355_out0[11:11];
assign v$_6815_out0 = v$CIN_2370_out0[11:11];
assign v$_7644_out0 = v$CIN_2355_out0[12:12];
assign v$_7659_out0 = v$CIN_2370_out0[12:12];
assign v$_8699_out0 = v$CIN_2355_out0[13:13];
assign v$_8714_out0 = v$CIN_2370_out0[13:13];
assign v$_8769_out0 = v$CIN_2355_out0[14:14];
assign v$_8784_out0 = v$CIN_2370_out0[14:14];
assign v$_10719_out0 = v$CIN_2355_out0[5:5];
assign v$_10734_out0 = v$CIN_2370_out0[5:5];
assign v$_13448_out0 = v$CIN_2355_out0[4:4];
assign v$_13463_out0 = v$CIN_2370_out0[4:4];
assign v$RM_3355_out0 = v$_7644_out0;
assign v$RM_3356_out0 = v$_8769_out0;
assign v$RM_3358_out0 = v$_10719_out0;
assign v$RM_3359_out0 = v$_13448_out0;
assign v$RM_3360_out0 = v$_8699_out0;
assign v$RM_3361_out0 = v$_3051_out0;
assign v$RM_3362_out0 = v$_3861_out0;
assign v$RM_3363_out0 = v$_3823_out0;
assign v$RM_3364_out0 = v$_2155_out0;
assign v$RM_3365_out0 = v$_1773_out0;
assign v$RM_3366_out0 = v$_3139_out0;
assign v$RM_3367_out0 = v$_6800_out0;
assign v$RM_3368_out0 = v$_468_out0;
assign v$RM_3369_out0 = v$_3085_out0;
assign v$RM_3579_out0 = v$_7659_out0;
assign v$RM_3580_out0 = v$_8784_out0;
assign v$RM_3582_out0 = v$_10734_out0;
assign v$RM_3583_out0 = v$_13463_out0;
assign v$RM_3584_out0 = v$_8714_out0;
assign v$RM_3585_out0 = v$_3066_out0;
assign v$RM_3586_out0 = v$_3876_out0;
assign v$RM_3587_out0 = v$_3838_out0;
assign v$RM_3588_out0 = v$_2170_out0;
assign v$RM_3589_out0 = v$_1788_out0;
assign v$RM_3590_out0 = v$_3154_out0;
assign v$RM_3591_out0 = v$_6815_out0;
assign v$RM_3592_out0 = v$_483_out0;
assign v$RM_3593_out0 = v$_3100_out0;
assign v$CIN_9810_out0 = v$_2195_out0;
assign v$CIN_10034_out0 = v$_2209_out0;
assign v$RM_11314_out0 = v$_2502_out0;
assign v$RM_11778_out0 = v$_2517_out0;
assign v$RD_5867_out0 = v$CIN_9810_out0;
assign v$RD_6331_out0 = v$CIN_10034_out0;
assign v$G1_7729_out0 = ((v$RD_5874_out0 && !v$RM_11314_out0) || (!v$RD_5874_out0) && v$RM_11314_out0);
assign v$G1_8193_out0 = ((v$RD_6338_out0 && !v$RM_11778_out0) || (!v$RD_6338_out0) && v$RM_11778_out0);
assign v$RM_11302_out0 = v$RM_3355_out0;
assign v$RM_11304_out0 = v$RM_3356_out0;
assign v$RM_11308_out0 = v$RM_3358_out0;
assign v$RM_11310_out0 = v$RM_3359_out0;
assign v$RM_11312_out0 = v$RM_3360_out0;
assign v$RM_11315_out0 = v$RM_3361_out0;
assign v$RM_11317_out0 = v$RM_3362_out0;
assign v$RM_11319_out0 = v$RM_3363_out0;
assign v$RM_11321_out0 = v$RM_3364_out0;
assign v$RM_11323_out0 = v$RM_3365_out0;
assign v$RM_11325_out0 = v$RM_3366_out0;
assign v$RM_11327_out0 = v$RM_3367_out0;
assign v$RM_11329_out0 = v$RM_3368_out0;
assign v$RM_11331_out0 = v$RM_3369_out0;
assign v$RM_11766_out0 = v$RM_3579_out0;
assign v$RM_11768_out0 = v$RM_3580_out0;
assign v$RM_11772_out0 = v$RM_3582_out0;
assign v$RM_11774_out0 = v$RM_3583_out0;
assign v$RM_11776_out0 = v$RM_3584_out0;
assign v$RM_11779_out0 = v$RM_3585_out0;
assign v$RM_11781_out0 = v$RM_3586_out0;
assign v$RM_11783_out0 = v$RM_3587_out0;
assign v$RM_11785_out0 = v$RM_3588_out0;
assign v$RM_11787_out0 = v$RM_3589_out0;
assign v$RM_11789_out0 = v$RM_3590_out0;
assign v$RM_11791_out0 = v$RM_3591_out0;
assign v$RM_11793_out0 = v$RM_3592_out0;
assign v$RM_11795_out0 = v$RM_3593_out0;
assign v$G2_12265_out0 = v$RD_5874_out0 && v$RM_11314_out0;
assign v$G2_12729_out0 = v$RD_6338_out0 && v$RM_11778_out0;
assign v$CARRY_4874_out0 = v$G2_12265_out0;
assign v$CARRY_5338_out0 = v$G2_12729_out0;
assign v$G1_7717_out0 = ((v$RD_5862_out0 && !v$RM_11302_out0) || (!v$RD_5862_out0) && v$RM_11302_out0);
assign v$G1_7719_out0 = ((v$RD_5864_out0 && !v$RM_11304_out0) || (!v$RD_5864_out0) && v$RM_11304_out0);
assign v$G1_7723_out0 = ((v$RD_5868_out0 && !v$RM_11308_out0) || (!v$RD_5868_out0) && v$RM_11308_out0);
assign v$G1_7725_out0 = ((v$RD_5870_out0 && !v$RM_11310_out0) || (!v$RD_5870_out0) && v$RM_11310_out0);
assign v$G1_7727_out0 = ((v$RD_5872_out0 && !v$RM_11312_out0) || (!v$RD_5872_out0) && v$RM_11312_out0);
assign v$G1_7730_out0 = ((v$RD_5875_out0 && !v$RM_11315_out0) || (!v$RD_5875_out0) && v$RM_11315_out0);
assign v$G1_7732_out0 = ((v$RD_5877_out0 && !v$RM_11317_out0) || (!v$RD_5877_out0) && v$RM_11317_out0);
assign v$G1_7734_out0 = ((v$RD_5879_out0 && !v$RM_11319_out0) || (!v$RD_5879_out0) && v$RM_11319_out0);
assign v$G1_7736_out0 = ((v$RD_5881_out0 && !v$RM_11321_out0) || (!v$RD_5881_out0) && v$RM_11321_out0);
assign v$G1_7738_out0 = ((v$RD_5883_out0 && !v$RM_11323_out0) || (!v$RD_5883_out0) && v$RM_11323_out0);
assign v$G1_7740_out0 = ((v$RD_5885_out0 && !v$RM_11325_out0) || (!v$RD_5885_out0) && v$RM_11325_out0);
assign v$G1_7742_out0 = ((v$RD_5887_out0 && !v$RM_11327_out0) || (!v$RD_5887_out0) && v$RM_11327_out0);
assign v$G1_7744_out0 = ((v$RD_5889_out0 && !v$RM_11329_out0) || (!v$RD_5889_out0) && v$RM_11329_out0);
assign v$G1_7746_out0 = ((v$RD_5891_out0 && !v$RM_11331_out0) || (!v$RD_5891_out0) && v$RM_11331_out0);
assign v$G1_8181_out0 = ((v$RD_6326_out0 && !v$RM_11766_out0) || (!v$RD_6326_out0) && v$RM_11766_out0);
assign v$G1_8183_out0 = ((v$RD_6328_out0 && !v$RM_11768_out0) || (!v$RD_6328_out0) && v$RM_11768_out0);
assign v$G1_8187_out0 = ((v$RD_6332_out0 && !v$RM_11772_out0) || (!v$RD_6332_out0) && v$RM_11772_out0);
assign v$G1_8189_out0 = ((v$RD_6334_out0 && !v$RM_11774_out0) || (!v$RD_6334_out0) && v$RM_11774_out0);
assign v$G1_8191_out0 = ((v$RD_6336_out0 && !v$RM_11776_out0) || (!v$RD_6336_out0) && v$RM_11776_out0);
assign v$G1_8194_out0 = ((v$RD_6339_out0 && !v$RM_11779_out0) || (!v$RD_6339_out0) && v$RM_11779_out0);
assign v$G1_8196_out0 = ((v$RD_6341_out0 && !v$RM_11781_out0) || (!v$RD_6341_out0) && v$RM_11781_out0);
assign v$G1_8198_out0 = ((v$RD_6343_out0 && !v$RM_11783_out0) || (!v$RD_6343_out0) && v$RM_11783_out0);
assign v$G1_8200_out0 = ((v$RD_6345_out0 && !v$RM_11785_out0) || (!v$RD_6345_out0) && v$RM_11785_out0);
assign v$G1_8202_out0 = ((v$RD_6347_out0 && !v$RM_11787_out0) || (!v$RD_6347_out0) && v$RM_11787_out0);
assign v$G1_8204_out0 = ((v$RD_6349_out0 && !v$RM_11789_out0) || (!v$RD_6349_out0) && v$RM_11789_out0);
assign v$G1_8206_out0 = ((v$RD_6351_out0 && !v$RM_11791_out0) || (!v$RD_6351_out0) && v$RM_11791_out0);
assign v$G1_8208_out0 = ((v$RD_6353_out0 && !v$RM_11793_out0) || (!v$RD_6353_out0) && v$RM_11793_out0);
assign v$G1_8210_out0 = ((v$RD_6355_out0 && !v$RM_11795_out0) || (!v$RD_6355_out0) && v$RM_11795_out0);
assign v$S_8875_out0 = v$G1_7729_out0;
assign v$S_9339_out0 = v$G1_8193_out0;
assign v$G2_12253_out0 = v$RD_5862_out0 && v$RM_11302_out0;
assign v$G2_12255_out0 = v$RD_5864_out0 && v$RM_11304_out0;
assign v$G2_12259_out0 = v$RD_5868_out0 && v$RM_11308_out0;
assign v$G2_12261_out0 = v$RD_5870_out0 && v$RM_11310_out0;
assign v$G2_12263_out0 = v$RD_5872_out0 && v$RM_11312_out0;
assign v$G2_12266_out0 = v$RD_5875_out0 && v$RM_11315_out0;
assign v$G2_12268_out0 = v$RD_5877_out0 && v$RM_11317_out0;
assign v$G2_12270_out0 = v$RD_5879_out0 && v$RM_11319_out0;
assign v$G2_12272_out0 = v$RD_5881_out0 && v$RM_11321_out0;
assign v$G2_12274_out0 = v$RD_5883_out0 && v$RM_11323_out0;
assign v$G2_12276_out0 = v$RD_5885_out0 && v$RM_11325_out0;
assign v$G2_12278_out0 = v$RD_5887_out0 && v$RM_11327_out0;
assign v$G2_12280_out0 = v$RD_5889_out0 && v$RM_11329_out0;
assign v$G2_12282_out0 = v$RD_5891_out0 && v$RM_11331_out0;
assign v$G2_12717_out0 = v$RD_6326_out0 && v$RM_11766_out0;
assign v$G2_12719_out0 = v$RD_6328_out0 && v$RM_11768_out0;
assign v$G2_12723_out0 = v$RD_6332_out0 && v$RM_11772_out0;
assign v$G2_12725_out0 = v$RD_6334_out0 && v$RM_11774_out0;
assign v$G2_12727_out0 = v$RD_6336_out0 && v$RM_11776_out0;
assign v$G2_12730_out0 = v$RD_6339_out0 && v$RM_11779_out0;
assign v$G2_12732_out0 = v$RD_6341_out0 && v$RM_11781_out0;
assign v$G2_12734_out0 = v$RD_6343_out0 && v$RM_11783_out0;
assign v$G2_12736_out0 = v$RD_6345_out0 && v$RM_11785_out0;
assign v$G2_12738_out0 = v$RD_6347_out0 && v$RM_11787_out0;
assign v$G2_12740_out0 = v$RD_6349_out0 && v$RM_11789_out0;
assign v$G2_12742_out0 = v$RD_6351_out0 && v$RM_11791_out0;
assign v$G2_12744_out0 = v$RD_6353_out0 && v$RM_11793_out0;
assign v$G2_12746_out0 = v$RD_6355_out0 && v$RM_11795_out0;
assign v$S_4665_out0 = v$S_8875_out0;
assign v$S_4680_out0 = v$S_9339_out0;
assign v$CARRY_4862_out0 = v$G2_12253_out0;
assign v$CARRY_4864_out0 = v$G2_12255_out0;
assign v$CARRY_4868_out0 = v$G2_12259_out0;
assign v$CARRY_4870_out0 = v$G2_12261_out0;
assign v$CARRY_4872_out0 = v$G2_12263_out0;
assign v$CARRY_4875_out0 = v$G2_12266_out0;
assign v$CARRY_4877_out0 = v$G2_12268_out0;
assign v$CARRY_4879_out0 = v$G2_12270_out0;
assign v$CARRY_4881_out0 = v$G2_12272_out0;
assign v$CARRY_4883_out0 = v$G2_12274_out0;
assign v$CARRY_4885_out0 = v$G2_12276_out0;
assign v$CARRY_4887_out0 = v$G2_12278_out0;
assign v$CARRY_4889_out0 = v$G2_12280_out0;
assign v$CARRY_4891_out0 = v$G2_12282_out0;
assign v$CARRY_5326_out0 = v$G2_12717_out0;
assign v$CARRY_5328_out0 = v$G2_12719_out0;
assign v$CARRY_5332_out0 = v$G2_12723_out0;
assign v$CARRY_5334_out0 = v$G2_12725_out0;
assign v$CARRY_5336_out0 = v$G2_12727_out0;
assign v$CARRY_5339_out0 = v$G2_12730_out0;
assign v$CARRY_5341_out0 = v$G2_12732_out0;
assign v$CARRY_5343_out0 = v$G2_12734_out0;
assign v$CARRY_5345_out0 = v$G2_12736_out0;
assign v$CARRY_5347_out0 = v$G2_12738_out0;
assign v$CARRY_5349_out0 = v$G2_12740_out0;
assign v$CARRY_5351_out0 = v$G2_12742_out0;
assign v$CARRY_5353_out0 = v$G2_12744_out0;
assign v$CARRY_5355_out0 = v$G2_12746_out0;
assign v$S_8863_out0 = v$G1_7717_out0;
assign v$S_8865_out0 = v$G1_7719_out0;
assign v$S_8869_out0 = v$G1_7723_out0;
assign v$S_8871_out0 = v$G1_7725_out0;
assign v$S_8873_out0 = v$G1_7727_out0;
assign v$S_8876_out0 = v$G1_7730_out0;
assign v$S_8878_out0 = v$G1_7732_out0;
assign v$S_8880_out0 = v$G1_7734_out0;
assign v$S_8882_out0 = v$G1_7736_out0;
assign v$S_8884_out0 = v$G1_7738_out0;
assign v$S_8886_out0 = v$G1_7740_out0;
assign v$S_8888_out0 = v$G1_7742_out0;
assign v$S_8890_out0 = v$G1_7744_out0;
assign v$S_8892_out0 = v$G1_7746_out0;
assign v$S_9327_out0 = v$G1_8181_out0;
assign v$S_9329_out0 = v$G1_8183_out0;
assign v$S_9333_out0 = v$G1_8187_out0;
assign v$S_9335_out0 = v$G1_8189_out0;
assign v$S_9337_out0 = v$G1_8191_out0;
assign v$S_9340_out0 = v$G1_8194_out0;
assign v$S_9342_out0 = v$G1_8196_out0;
assign v$S_9344_out0 = v$G1_8198_out0;
assign v$S_9346_out0 = v$G1_8200_out0;
assign v$S_9348_out0 = v$G1_8202_out0;
assign v$S_9350_out0 = v$G1_8204_out0;
assign v$S_9352_out0 = v$G1_8206_out0;
assign v$S_9354_out0 = v$G1_8208_out0;
assign v$S_9356_out0 = v$G1_8210_out0;
assign v$CIN_9816_out0 = v$CARRY_4874_out0;
assign v$CIN_10040_out0 = v$CARRY_5338_out0;
assign v$_2392_out0 = { v$_4529_out0,v$S_4665_out0 };
assign v$_2393_out0 = { v$_4530_out0,v$S_4680_out0 };
assign v$RD_5880_out0 = v$CIN_9816_out0;
assign v$RD_6344_out0 = v$CIN_10040_out0;
assign v$RM_11303_out0 = v$S_8863_out0;
assign v$RM_11305_out0 = v$S_8865_out0;
assign v$RM_11309_out0 = v$S_8869_out0;
assign v$RM_11311_out0 = v$S_8871_out0;
assign v$RM_11313_out0 = v$S_8873_out0;
assign v$RM_11316_out0 = v$S_8876_out0;
assign v$RM_11318_out0 = v$S_8878_out0;
assign v$RM_11320_out0 = v$S_8880_out0;
assign v$RM_11322_out0 = v$S_8882_out0;
assign v$RM_11324_out0 = v$S_8884_out0;
assign v$RM_11326_out0 = v$S_8886_out0;
assign v$RM_11328_out0 = v$S_8888_out0;
assign v$RM_11330_out0 = v$S_8890_out0;
assign v$RM_11332_out0 = v$S_8892_out0;
assign v$RM_11767_out0 = v$S_9327_out0;
assign v$RM_11769_out0 = v$S_9329_out0;
assign v$RM_11773_out0 = v$S_9333_out0;
assign v$RM_11775_out0 = v$S_9335_out0;
assign v$RM_11777_out0 = v$S_9337_out0;
assign v$RM_11780_out0 = v$S_9340_out0;
assign v$RM_11782_out0 = v$S_9342_out0;
assign v$RM_11784_out0 = v$S_9344_out0;
assign v$RM_11786_out0 = v$S_9346_out0;
assign v$RM_11788_out0 = v$S_9348_out0;
assign v$RM_11790_out0 = v$S_9350_out0;
assign v$RM_11792_out0 = v$S_9352_out0;
assign v$RM_11794_out0 = v$S_9354_out0;
assign v$RM_11796_out0 = v$S_9356_out0;
assign v$G1_7735_out0 = ((v$RD_5880_out0 && !v$RM_11320_out0) || (!v$RD_5880_out0) && v$RM_11320_out0);
assign v$G1_8199_out0 = ((v$RD_6344_out0 && !v$RM_11784_out0) || (!v$RD_6344_out0) && v$RM_11784_out0);
assign v$G2_12271_out0 = v$RD_5880_out0 && v$RM_11320_out0;
assign v$G2_12735_out0 = v$RD_6344_out0 && v$RM_11784_out0;
assign v$CARRY_4880_out0 = v$G2_12271_out0;
assign v$CARRY_5344_out0 = v$G2_12735_out0;
assign v$S_8881_out0 = v$G1_7735_out0;
assign v$S_9345_out0 = v$G1_8199_out0;
assign v$S_1227_out0 = v$S_8881_out0;
assign v$S_1451_out0 = v$S_9345_out0;
assign v$G1_4003_out0 = v$CARRY_4880_out0 || v$CARRY_4879_out0;
assign v$G1_4227_out0 = v$CARRY_5344_out0 || v$CARRY_5343_out0;
assign v$COUT_695_out0 = v$G1_4003_out0;
assign v$COUT_919_out0 = v$G1_4227_out0;
assign v$CIN_9822_out0 = v$COUT_695_out0;
assign v$CIN_10046_out0 = v$COUT_919_out0;
assign v$RD_5892_out0 = v$CIN_9822_out0;
assign v$RD_6356_out0 = v$CIN_10046_out0;
assign v$G1_7747_out0 = ((v$RD_5892_out0 && !v$RM_11332_out0) || (!v$RD_5892_out0) && v$RM_11332_out0);
assign v$G1_8211_out0 = ((v$RD_6356_out0 && !v$RM_11796_out0) || (!v$RD_6356_out0) && v$RM_11796_out0);
assign v$G2_12283_out0 = v$RD_5892_out0 && v$RM_11332_out0;
assign v$G2_12747_out0 = v$RD_6356_out0 && v$RM_11796_out0;
assign v$CARRY_4892_out0 = v$G2_12283_out0;
assign v$CARRY_5356_out0 = v$G2_12747_out0;
assign v$S_8893_out0 = v$G1_7747_out0;
assign v$S_9357_out0 = v$G1_8211_out0;
assign v$S_1233_out0 = v$S_8893_out0;
assign v$S_1457_out0 = v$S_9357_out0;
assign v$G1_4009_out0 = v$CARRY_4892_out0 || v$CARRY_4891_out0;
assign v$G1_4233_out0 = v$CARRY_5356_out0 || v$CARRY_5355_out0;
assign v$COUT_701_out0 = v$G1_4009_out0;
assign v$COUT_925_out0 = v$G1_4233_out0;
assign v$_4782_out0 = { v$S_1227_out0,v$S_1233_out0 };
assign v$_4797_out0 = { v$S_1451_out0,v$S_1457_out0 };
assign v$CIN_9817_out0 = v$COUT_701_out0;
assign v$CIN_10041_out0 = v$COUT_925_out0;
assign v$RD_5882_out0 = v$CIN_9817_out0;
assign v$RD_6346_out0 = v$CIN_10041_out0;
assign v$G1_7737_out0 = ((v$RD_5882_out0 && !v$RM_11322_out0) || (!v$RD_5882_out0) && v$RM_11322_out0);
assign v$G1_8201_out0 = ((v$RD_6346_out0 && !v$RM_11786_out0) || (!v$RD_6346_out0) && v$RM_11786_out0);
assign v$G2_12273_out0 = v$RD_5882_out0 && v$RM_11322_out0;
assign v$G2_12737_out0 = v$RD_6346_out0 && v$RM_11786_out0;
assign v$CARRY_4882_out0 = v$G2_12273_out0;
assign v$CARRY_5346_out0 = v$G2_12737_out0;
assign v$S_8883_out0 = v$G1_7737_out0;
assign v$S_9347_out0 = v$G1_8201_out0;
assign v$S_1228_out0 = v$S_8883_out0;
assign v$S_1452_out0 = v$S_9347_out0;
assign v$G1_4004_out0 = v$CARRY_4882_out0 || v$CARRY_4881_out0;
assign v$G1_4228_out0 = v$CARRY_5346_out0 || v$CARRY_5345_out0;
assign v$COUT_696_out0 = v$G1_4004_out0;
assign v$COUT_920_out0 = v$G1_4228_out0;
assign v$_2552_out0 = { v$_4782_out0,v$S_1228_out0 };
assign v$_2567_out0 = { v$_4797_out0,v$S_1452_out0 };
assign v$CIN_9812_out0 = v$COUT_696_out0;
assign v$CIN_10036_out0 = v$COUT_920_out0;
assign v$RD_5871_out0 = v$CIN_9812_out0;
assign v$RD_6335_out0 = v$CIN_10036_out0;
assign v$G1_7726_out0 = ((v$RD_5871_out0 && !v$RM_11311_out0) || (!v$RD_5871_out0) && v$RM_11311_out0);
assign v$G1_8190_out0 = ((v$RD_6335_out0 && !v$RM_11775_out0) || (!v$RD_6335_out0) && v$RM_11775_out0);
assign v$G2_12262_out0 = v$RD_5871_out0 && v$RM_11311_out0;
assign v$G2_12726_out0 = v$RD_6335_out0 && v$RM_11775_out0;
assign v$CARRY_4871_out0 = v$G2_12262_out0;
assign v$CARRY_5335_out0 = v$G2_12726_out0;
assign v$S_8872_out0 = v$G1_7726_out0;
assign v$S_9336_out0 = v$G1_8190_out0;
assign v$S_1223_out0 = v$S_8872_out0;
assign v$S_1447_out0 = v$S_9336_out0;
assign v$G1_3999_out0 = v$CARRY_4871_out0 || v$CARRY_4870_out0;
assign v$G1_4223_out0 = v$CARRY_5335_out0 || v$CARRY_5334_out0;
assign v$COUT_691_out0 = v$G1_3999_out0;
assign v$COUT_915_out0 = v$G1_4223_out0;
assign v$_7032_out0 = { v$_2552_out0,v$S_1223_out0 };
assign v$_7047_out0 = { v$_2567_out0,v$S_1447_out0 };
assign v$CIN_9811_out0 = v$COUT_691_out0;
assign v$CIN_10035_out0 = v$COUT_915_out0;
assign v$RD_5869_out0 = v$CIN_9811_out0;
assign v$RD_6333_out0 = v$CIN_10035_out0;
assign v$G1_7724_out0 = ((v$RD_5869_out0 && !v$RM_11309_out0) || (!v$RD_5869_out0) && v$RM_11309_out0);
assign v$G1_8188_out0 = ((v$RD_6333_out0 && !v$RM_11773_out0) || (!v$RD_6333_out0) && v$RM_11773_out0);
assign v$G2_12260_out0 = v$RD_5869_out0 && v$RM_11309_out0;
assign v$G2_12724_out0 = v$RD_6333_out0 && v$RM_11773_out0;
assign v$CARRY_4869_out0 = v$G2_12260_out0;
assign v$CARRY_5333_out0 = v$G2_12724_out0;
assign v$S_8870_out0 = v$G1_7724_out0;
assign v$S_9334_out0 = v$G1_8188_out0;
assign v$S_1222_out0 = v$S_8870_out0;
assign v$S_1446_out0 = v$S_9334_out0;
assign v$G1_3998_out0 = v$CARRY_4869_out0 || v$CARRY_4868_out0;
assign v$G1_4222_out0 = v$CARRY_5333_out0 || v$CARRY_5332_out0;
assign v$COUT_690_out0 = v$G1_3998_out0;
assign v$COUT_914_out0 = v$G1_4222_out0;
assign v$_13518_out0 = { v$_7032_out0,v$S_1222_out0 };
assign v$_13533_out0 = { v$_7047_out0,v$S_1446_out0 };
assign v$CIN_9818_out0 = v$COUT_690_out0;
assign v$CIN_10042_out0 = v$COUT_914_out0;
assign v$RD_5884_out0 = v$CIN_9818_out0;
assign v$RD_6348_out0 = v$CIN_10042_out0;
assign v$G1_7739_out0 = ((v$RD_5884_out0 && !v$RM_11324_out0) || (!v$RD_5884_out0) && v$RM_11324_out0);
assign v$G1_8203_out0 = ((v$RD_6348_out0 && !v$RM_11788_out0) || (!v$RD_6348_out0) && v$RM_11788_out0);
assign v$G2_12275_out0 = v$RD_5884_out0 && v$RM_11324_out0;
assign v$G2_12739_out0 = v$RD_6348_out0 && v$RM_11788_out0;
assign v$CARRY_4884_out0 = v$G2_12275_out0;
assign v$CARRY_5348_out0 = v$G2_12739_out0;
assign v$S_8885_out0 = v$G1_7739_out0;
assign v$S_9349_out0 = v$G1_8203_out0;
assign v$S_1229_out0 = v$S_8885_out0;
assign v$S_1453_out0 = v$S_9349_out0;
assign v$G1_4005_out0 = v$CARRY_4884_out0 || v$CARRY_4883_out0;
assign v$G1_4229_out0 = v$CARRY_5348_out0 || v$CARRY_5347_out0;
assign v$COUT_697_out0 = v$G1_4005_out0;
assign v$COUT_921_out0 = v$G1_4229_out0;
assign v$_3311_out0 = { v$_13518_out0,v$S_1229_out0 };
assign v$_3326_out0 = { v$_13533_out0,v$S_1453_out0 };
assign v$CIN_9819_out0 = v$COUT_697_out0;
assign v$CIN_10043_out0 = v$COUT_921_out0;
assign v$RD_5886_out0 = v$CIN_9819_out0;
assign v$RD_6350_out0 = v$CIN_10043_out0;
assign v$G1_7741_out0 = ((v$RD_5886_out0 && !v$RM_11326_out0) || (!v$RD_5886_out0) && v$RM_11326_out0);
assign v$G1_8205_out0 = ((v$RD_6350_out0 && !v$RM_11790_out0) || (!v$RD_6350_out0) && v$RM_11790_out0);
assign v$G2_12277_out0 = v$RD_5886_out0 && v$RM_11326_out0;
assign v$G2_12741_out0 = v$RD_6350_out0 && v$RM_11790_out0;
assign v$CARRY_4886_out0 = v$G2_12277_out0;
assign v$CARRY_5350_out0 = v$G2_12741_out0;
assign v$S_8887_out0 = v$G1_7741_out0;
assign v$S_9351_out0 = v$G1_8205_out0;
assign v$S_1230_out0 = v$S_8887_out0;
assign v$S_1454_out0 = v$S_9351_out0;
assign v$G1_4006_out0 = v$CARRY_4886_out0 || v$CARRY_4885_out0;
assign v$G1_4230_out0 = v$CARRY_5350_out0 || v$CARRY_5349_out0;
assign v$COUT_698_out0 = v$G1_4006_out0;
assign v$COUT_922_out0 = v$G1_4230_out0;
assign v$_7147_out0 = { v$_3311_out0,v$S_1230_out0 };
assign v$_7162_out0 = { v$_3326_out0,v$S_1454_out0 };
assign v$CIN_9821_out0 = v$COUT_698_out0;
assign v$CIN_10045_out0 = v$COUT_922_out0;
assign v$RD_5890_out0 = v$CIN_9821_out0;
assign v$RD_6354_out0 = v$CIN_10045_out0;
assign v$G1_7745_out0 = ((v$RD_5890_out0 && !v$RM_11330_out0) || (!v$RD_5890_out0) && v$RM_11330_out0);
assign v$G1_8209_out0 = ((v$RD_6354_out0 && !v$RM_11794_out0) || (!v$RD_6354_out0) && v$RM_11794_out0);
assign v$G2_12281_out0 = v$RD_5890_out0 && v$RM_11330_out0;
assign v$G2_12745_out0 = v$RD_6354_out0 && v$RM_11794_out0;
assign v$CARRY_4890_out0 = v$G2_12281_out0;
assign v$CARRY_5354_out0 = v$G2_12745_out0;
assign v$S_8891_out0 = v$G1_7745_out0;
assign v$S_9355_out0 = v$G1_8209_out0;
assign v$S_1232_out0 = v$S_8891_out0;
assign v$S_1456_out0 = v$S_9355_out0;
assign v$G1_4008_out0 = v$CARRY_4890_out0 || v$CARRY_4889_out0;
assign v$G1_4232_out0 = v$CARRY_5354_out0 || v$CARRY_5353_out0;
assign v$COUT_700_out0 = v$G1_4008_out0;
assign v$COUT_924_out0 = v$G1_4232_out0;
assign v$_4749_out0 = { v$_7147_out0,v$S_1232_out0 };
assign v$_4764_out0 = { v$_7162_out0,v$S_1456_out0 };
assign v$CIN_9814_out0 = v$COUT_700_out0;
assign v$CIN_10038_out0 = v$COUT_924_out0;
assign v$RD_5876_out0 = v$CIN_9814_out0;
assign v$RD_6340_out0 = v$CIN_10038_out0;
assign v$G1_7731_out0 = ((v$RD_5876_out0 && !v$RM_11316_out0) || (!v$RD_5876_out0) && v$RM_11316_out0);
assign v$G1_8195_out0 = ((v$RD_6340_out0 && !v$RM_11780_out0) || (!v$RD_6340_out0) && v$RM_11780_out0);
assign v$G2_12267_out0 = v$RD_5876_out0 && v$RM_11316_out0;
assign v$G2_12731_out0 = v$RD_6340_out0 && v$RM_11780_out0;
assign v$CARRY_4876_out0 = v$G2_12267_out0;
assign v$CARRY_5340_out0 = v$G2_12731_out0;
assign v$S_8877_out0 = v$G1_7731_out0;
assign v$S_9341_out0 = v$G1_8195_out0;
assign v$S_1225_out0 = v$S_8877_out0;
assign v$S_1449_out0 = v$S_9341_out0;
assign v$G1_4001_out0 = v$CARRY_4876_out0 || v$CARRY_4875_out0;
assign v$G1_4225_out0 = v$CARRY_5340_out0 || v$CARRY_5339_out0;
assign v$COUT_693_out0 = v$G1_4001_out0;
assign v$COUT_917_out0 = v$G1_4225_out0;
assign v$_6926_out0 = { v$_4749_out0,v$S_1225_out0 };
assign v$_6941_out0 = { v$_4764_out0,v$S_1449_out0 };
assign v$CIN_9815_out0 = v$COUT_693_out0;
assign v$CIN_10039_out0 = v$COUT_917_out0;
assign v$RD_5878_out0 = v$CIN_9815_out0;
assign v$RD_6342_out0 = v$CIN_10039_out0;
assign v$G1_7733_out0 = ((v$RD_5878_out0 && !v$RM_11318_out0) || (!v$RD_5878_out0) && v$RM_11318_out0);
assign v$G1_8197_out0 = ((v$RD_6342_out0 && !v$RM_11782_out0) || (!v$RD_6342_out0) && v$RM_11782_out0);
assign v$G2_12269_out0 = v$RD_5878_out0 && v$RM_11318_out0;
assign v$G2_12733_out0 = v$RD_6342_out0 && v$RM_11782_out0;
assign v$CARRY_4878_out0 = v$G2_12269_out0;
assign v$CARRY_5342_out0 = v$G2_12733_out0;
assign v$S_8879_out0 = v$G1_7733_out0;
assign v$S_9343_out0 = v$G1_8197_out0;
assign v$S_1226_out0 = v$S_8879_out0;
assign v$S_1450_out0 = v$S_9343_out0;
assign v$G1_4002_out0 = v$CARRY_4878_out0 || v$CARRY_4877_out0;
assign v$G1_4226_out0 = v$CARRY_5342_out0 || v$CARRY_5341_out0;
assign v$COUT_694_out0 = v$G1_4002_out0;
assign v$COUT_918_out0 = v$G1_4226_out0;
assign v$_5802_out0 = { v$_6926_out0,v$S_1226_out0 };
assign v$_5817_out0 = { v$_6941_out0,v$S_1450_out0 };
assign v$CIN_9820_out0 = v$COUT_694_out0;
assign v$CIN_10044_out0 = v$COUT_918_out0;
assign v$RD_5888_out0 = v$CIN_9820_out0;
assign v$RD_6352_out0 = v$CIN_10044_out0;
assign v$G1_7743_out0 = ((v$RD_5888_out0 && !v$RM_11328_out0) || (!v$RD_5888_out0) && v$RM_11328_out0);
assign v$G1_8207_out0 = ((v$RD_6352_out0 && !v$RM_11792_out0) || (!v$RD_6352_out0) && v$RM_11792_out0);
assign v$G2_12279_out0 = v$RD_5888_out0 && v$RM_11328_out0;
assign v$G2_12743_out0 = v$RD_6352_out0 && v$RM_11792_out0;
assign v$CARRY_4888_out0 = v$G2_12279_out0;
assign v$CARRY_5352_out0 = v$G2_12743_out0;
assign v$S_8889_out0 = v$G1_7743_out0;
assign v$S_9353_out0 = v$G1_8207_out0;
assign v$S_1231_out0 = v$S_8889_out0;
assign v$S_1455_out0 = v$S_9353_out0;
assign v$G1_4007_out0 = v$CARRY_4888_out0 || v$CARRY_4887_out0;
assign v$G1_4231_out0 = v$CARRY_5352_out0 || v$CARRY_5351_out0;
assign v$COUT_699_out0 = v$G1_4007_out0;
assign v$COUT_923_out0 = v$G1_4231_out0;
assign v$_2026_out0 = { v$_5802_out0,v$S_1231_out0 };
assign v$_2041_out0 = { v$_5817_out0,v$S_1455_out0 };
assign v$CIN_9808_out0 = v$COUT_699_out0;
assign v$CIN_10032_out0 = v$COUT_923_out0;
assign v$RD_5863_out0 = v$CIN_9808_out0;
assign v$RD_6327_out0 = v$CIN_10032_out0;
assign v$G1_7718_out0 = ((v$RD_5863_out0 && !v$RM_11303_out0) || (!v$RD_5863_out0) && v$RM_11303_out0);
assign v$G1_8182_out0 = ((v$RD_6327_out0 && !v$RM_11767_out0) || (!v$RD_6327_out0) && v$RM_11767_out0);
assign v$G2_12254_out0 = v$RD_5863_out0 && v$RM_11303_out0;
assign v$G2_12718_out0 = v$RD_6327_out0 && v$RM_11767_out0;
assign v$CARRY_4863_out0 = v$G2_12254_out0;
assign v$CARRY_5327_out0 = v$G2_12718_out0;
assign v$S_8864_out0 = v$G1_7718_out0;
assign v$S_9328_out0 = v$G1_8182_out0;
assign v$S_1219_out0 = v$S_8864_out0;
assign v$S_1443_out0 = v$S_9328_out0;
assign v$G1_3995_out0 = v$CARRY_4863_out0 || v$CARRY_4862_out0;
assign v$G1_4219_out0 = v$CARRY_5327_out0 || v$CARRY_5326_out0;
assign v$COUT_687_out0 = v$G1_3995_out0;
assign v$COUT_911_out0 = v$G1_4219_out0;
assign v$_2793_out0 = { v$_2026_out0,v$S_1219_out0 };
assign v$_2808_out0 = { v$_2041_out0,v$S_1443_out0 };
assign v$CIN_9813_out0 = v$COUT_687_out0;
assign v$CIN_10037_out0 = v$COUT_911_out0;
assign v$RD_5873_out0 = v$CIN_9813_out0;
assign v$RD_6337_out0 = v$CIN_10037_out0;
assign v$G1_7728_out0 = ((v$RD_5873_out0 && !v$RM_11313_out0) || (!v$RD_5873_out0) && v$RM_11313_out0);
assign v$G1_8192_out0 = ((v$RD_6337_out0 && !v$RM_11777_out0) || (!v$RD_6337_out0) && v$RM_11777_out0);
assign v$G2_12264_out0 = v$RD_5873_out0 && v$RM_11313_out0;
assign v$G2_12728_out0 = v$RD_6337_out0 && v$RM_11777_out0;
assign v$CARRY_4873_out0 = v$G2_12264_out0;
assign v$CARRY_5337_out0 = v$G2_12728_out0;
assign v$S_8874_out0 = v$G1_7728_out0;
assign v$S_9338_out0 = v$G1_8192_out0;
assign v$S_1224_out0 = v$S_8874_out0;
assign v$S_1448_out0 = v$S_9338_out0;
assign v$G1_4000_out0 = v$CARRY_4873_out0 || v$CARRY_4872_out0;
assign v$G1_4224_out0 = v$CARRY_5337_out0 || v$CARRY_5336_out0;
assign v$COUT_692_out0 = v$G1_4000_out0;
assign v$COUT_916_out0 = v$G1_4224_out0;
assign v$_1825_out0 = { v$_2793_out0,v$S_1224_out0 };
assign v$_1840_out0 = { v$_2808_out0,v$S_1448_out0 };
assign v$CIN_9809_out0 = v$COUT_692_out0;
assign v$CIN_10033_out0 = v$COUT_916_out0;
assign v$RD_5865_out0 = v$CIN_9809_out0;
assign v$RD_6329_out0 = v$CIN_10033_out0;
assign v$G1_7720_out0 = ((v$RD_5865_out0 && !v$RM_11305_out0) || (!v$RD_5865_out0) && v$RM_11305_out0);
assign v$G1_8184_out0 = ((v$RD_6329_out0 && !v$RM_11769_out0) || (!v$RD_6329_out0) && v$RM_11769_out0);
assign v$G2_12256_out0 = v$RD_5865_out0 && v$RM_11305_out0;
assign v$G2_12720_out0 = v$RD_6329_out0 && v$RM_11769_out0;
assign v$CARRY_4865_out0 = v$G2_12256_out0;
assign v$CARRY_5329_out0 = v$G2_12720_out0;
assign v$S_8866_out0 = v$G1_7720_out0;
assign v$S_9330_out0 = v$G1_8184_out0;
assign v$S_1220_out0 = v$S_8866_out0;
assign v$S_1444_out0 = v$S_9330_out0;
assign v$G1_3996_out0 = v$CARRY_4865_out0 || v$CARRY_4864_out0;
assign v$G1_4220_out0 = v$CARRY_5329_out0 || v$CARRY_5328_out0;
assign v$COUT_688_out0 = v$G1_3996_out0;
assign v$COUT_912_out0 = v$G1_4220_out0;
assign v$_4549_out0 = { v$_1825_out0,v$S_1220_out0 };
assign v$_4564_out0 = { v$_1840_out0,v$S_1444_out0 };
assign v$RM_3357_out0 = v$COUT_688_out0;
assign v$RM_3581_out0 = v$COUT_912_out0;
assign v$RM_11306_out0 = v$RM_3357_out0;
assign v$RM_11770_out0 = v$RM_3581_out0;
assign v$G1_7721_out0 = ((v$RD_5866_out0 && !v$RM_11306_out0) || (!v$RD_5866_out0) && v$RM_11306_out0);
assign v$G1_8185_out0 = ((v$RD_6330_out0 && !v$RM_11770_out0) || (!v$RD_6330_out0) && v$RM_11770_out0);
assign v$G2_12257_out0 = v$RD_5866_out0 && v$RM_11306_out0;
assign v$G2_12721_out0 = v$RD_6330_out0 && v$RM_11770_out0;
assign v$CARRY_4866_out0 = v$G2_12257_out0;
assign v$CARRY_5330_out0 = v$G2_12721_out0;
assign v$S_8867_out0 = v$G1_7721_out0;
assign v$S_9331_out0 = v$G1_8185_out0;
assign v$RM_11307_out0 = v$S_8867_out0;
assign v$RM_11771_out0 = v$S_9331_out0;
assign v$G1_7722_out0 = ((v$RD_5867_out0 && !v$RM_11307_out0) || (!v$RD_5867_out0) && v$RM_11307_out0);
assign v$G1_8186_out0 = ((v$RD_6331_out0 && !v$RM_11771_out0) || (!v$RD_6331_out0) && v$RM_11771_out0);
assign v$G2_12258_out0 = v$RD_5867_out0 && v$RM_11307_out0;
assign v$G2_12722_out0 = v$RD_6331_out0 && v$RM_11771_out0;
assign v$CARRY_4867_out0 = v$G2_12258_out0;
assign v$CARRY_5331_out0 = v$G2_12722_out0;
assign v$S_8868_out0 = v$G1_7722_out0;
assign v$S_9332_out0 = v$G1_8186_out0;
assign v$S_1221_out0 = v$S_8868_out0;
assign v$S_1445_out0 = v$S_9332_out0;
assign v$G1_3997_out0 = v$CARRY_4867_out0 || v$CARRY_4866_out0;
assign v$G1_4221_out0 = v$CARRY_5331_out0 || v$CARRY_5330_out0;
assign v$COUT_689_out0 = v$G1_3997_out0;
assign v$COUT_913_out0 = v$G1_4221_out0;
assign v$_10651_out0 = { v$_4549_out0,v$S_1221_out0 };
assign v$_10666_out0 = { v$_4564_out0,v$S_1445_out0 };
assign v$_10946_out0 = { v$_10651_out0,v$COUT_689_out0 };
assign v$_10961_out0 = { v$_10666_out0,v$COUT_913_out0 };
assign v$COUT_10916_out0 = v$_10946_out0;
assign v$COUT_10931_out0 = v$_10961_out0;
assign v$CIN_2365_out0 = v$COUT_10916_out0;
assign v$CIN_2380_out0 = v$COUT_10931_out0;
assign v$_478_out0 = v$CIN_2365_out0[8:8];
assign v$_493_out0 = v$CIN_2380_out0[8:8];
assign v$_1783_out0 = v$CIN_2365_out0[6:6];
assign v$_1798_out0 = v$CIN_2380_out0[6:6];
assign v$_2165_out0 = v$CIN_2365_out0[3:3];
assign v$_2180_out0 = v$CIN_2380_out0[3:3];
assign v$_2204_out0 = v$CIN_2365_out0[15:15];
assign v$_2218_out0 = v$CIN_2380_out0[15:15];
assign v$_2512_out0 = v$CIN_2365_out0[0:0];
assign v$_2527_out0 = v$CIN_2380_out0[0:0];
assign v$_3061_out0 = v$CIN_2365_out0[9:9];
assign v$_3076_out0 = v$CIN_2380_out0[9:9];
assign v$_3095_out0 = v$CIN_2365_out0[2:2];
assign v$_3110_out0 = v$CIN_2380_out0[2:2];
assign v$_3149_out0 = v$CIN_2365_out0[7:7];
assign v$_3164_out0 = v$CIN_2380_out0[7:7];
assign v$_3833_out0 = v$CIN_2365_out0[1:1];
assign v$_3848_out0 = v$CIN_2380_out0[1:1];
assign v$_3871_out0 = v$CIN_2365_out0[10:10];
assign v$_3886_out0 = v$CIN_2380_out0[10:10];
assign v$_6810_out0 = v$CIN_2365_out0[11:11];
assign v$_6825_out0 = v$CIN_2380_out0[11:11];
assign v$_7654_out0 = v$CIN_2365_out0[12:12];
assign v$_7669_out0 = v$CIN_2380_out0[12:12];
assign v$_8709_out0 = v$CIN_2365_out0[13:13];
assign v$_8724_out0 = v$CIN_2380_out0[13:13];
assign v$_8779_out0 = v$CIN_2365_out0[14:14];
assign v$_8794_out0 = v$CIN_2380_out0[14:14];
assign v$_10729_out0 = v$CIN_2365_out0[5:5];
assign v$_10744_out0 = v$CIN_2380_out0[5:5];
assign v$_13458_out0 = v$CIN_2365_out0[4:4];
assign v$_13473_out0 = v$CIN_2380_out0[4:4];
assign v$RM_3504_out0 = v$_7654_out0;
assign v$RM_3505_out0 = v$_8779_out0;
assign v$RM_3507_out0 = v$_10729_out0;
assign v$RM_3508_out0 = v$_13458_out0;
assign v$RM_3509_out0 = v$_8709_out0;
assign v$RM_3510_out0 = v$_3061_out0;
assign v$RM_3511_out0 = v$_3871_out0;
assign v$RM_3512_out0 = v$_3833_out0;
assign v$RM_3513_out0 = v$_2165_out0;
assign v$RM_3514_out0 = v$_1783_out0;
assign v$RM_3515_out0 = v$_3149_out0;
assign v$RM_3516_out0 = v$_6810_out0;
assign v$RM_3517_out0 = v$_478_out0;
assign v$RM_3518_out0 = v$_3095_out0;
assign v$RM_3728_out0 = v$_7669_out0;
assign v$RM_3729_out0 = v$_8794_out0;
assign v$RM_3731_out0 = v$_10744_out0;
assign v$RM_3732_out0 = v$_13473_out0;
assign v$RM_3733_out0 = v$_8724_out0;
assign v$RM_3734_out0 = v$_3076_out0;
assign v$RM_3735_out0 = v$_3886_out0;
assign v$RM_3736_out0 = v$_3848_out0;
assign v$RM_3737_out0 = v$_2180_out0;
assign v$RM_3738_out0 = v$_1798_out0;
assign v$RM_3739_out0 = v$_3164_out0;
assign v$RM_3740_out0 = v$_6825_out0;
assign v$RM_3741_out0 = v$_493_out0;
assign v$RM_3742_out0 = v$_3110_out0;
assign v$CIN_9959_out0 = v$_2204_out0;
assign v$CIN_10183_out0 = v$_2218_out0;
assign v$RM_11623_out0 = v$_2512_out0;
assign v$RM_12087_out0 = v$_2527_out0;
assign v$RD_6176_out0 = v$CIN_9959_out0;
assign v$RD_6640_out0 = v$CIN_10183_out0;
assign v$G1_8038_out0 = ((v$RD_6183_out0 && !v$RM_11623_out0) || (!v$RD_6183_out0) && v$RM_11623_out0);
assign v$G1_8502_out0 = ((v$RD_6647_out0 && !v$RM_12087_out0) || (!v$RD_6647_out0) && v$RM_12087_out0);
assign v$RM_11611_out0 = v$RM_3504_out0;
assign v$RM_11613_out0 = v$RM_3505_out0;
assign v$RM_11617_out0 = v$RM_3507_out0;
assign v$RM_11619_out0 = v$RM_3508_out0;
assign v$RM_11621_out0 = v$RM_3509_out0;
assign v$RM_11624_out0 = v$RM_3510_out0;
assign v$RM_11626_out0 = v$RM_3511_out0;
assign v$RM_11628_out0 = v$RM_3512_out0;
assign v$RM_11630_out0 = v$RM_3513_out0;
assign v$RM_11632_out0 = v$RM_3514_out0;
assign v$RM_11634_out0 = v$RM_3515_out0;
assign v$RM_11636_out0 = v$RM_3516_out0;
assign v$RM_11638_out0 = v$RM_3517_out0;
assign v$RM_11640_out0 = v$RM_3518_out0;
assign v$RM_12075_out0 = v$RM_3728_out0;
assign v$RM_12077_out0 = v$RM_3729_out0;
assign v$RM_12081_out0 = v$RM_3731_out0;
assign v$RM_12083_out0 = v$RM_3732_out0;
assign v$RM_12085_out0 = v$RM_3733_out0;
assign v$RM_12088_out0 = v$RM_3734_out0;
assign v$RM_12090_out0 = v$RM_3735_out0;
assign v$RM_12092_out0 = v$RM_3736_out0;
assign v$RM_12094_out0 = v$RM_3737_out0;
assign v$RM_12096_out0 = v$RM_3738_out0;
assign v$RM_12098_out0 = v$RM_3739_out0;
assign v$RM_12100_out0 = v$RM_3740_out0;
assign v$RM_12102_out0 = v$RM_3741_out0;
assign v$RM_12104_out0 = v$RM_3742_out0;
assign v$G2_12574_out0 = v$RD_6183_out0 && v$RM_11623_out0;
assign v$G2_13038_out0 = v$RD_6647_out0 && v$RM_12087_out0;
assign v$CARRY_5183_out0 = v$G2_12574_out0;
assign v$CARRY_5647_out0 = v$G2_13038_out0;
assign v$G1_8026_out0 = ((v$RD_6171_out0 && !v$RM_11611_out0) || (!v$RD_6171_out0) && v$RM_11611_out0);
assign v$G1_8028_out0 = ((v$RD_6173_out0 && !v$RM_11613_out0) || (!v$RD_6173_out0) && v$RM_11613_out0);
assign v$G1_8032_out0 = ((v$RD_6177_out0 && !v$RM_11617_out0) || (!v$RD_6177_out0) && v$RM_11617_out0);
assign v$G1_8034_out0 = ((v$RD_6179_out0 && !v$RM_11619_out0) || (!v$RD_6179_out0) && v$RM_11619_out0);
assign v$G1_8036_out0 = ((v$RD_6181_out0 && !v$RM_11621_out0) || (!v$RD_6181_out0) && v$RM_11621_out0);
assign v$G1_8039_out0 = ((v$RD_6184_out0 && !v$RM_11624_out0) || (!v$RD_6184_out0) && v$RM_11624_out0);
assign v$G1_8041_out0 = ((v$RD_6186_out0 && !v$RM_11626_out0) || (!v$RD_6186_out0) && v$RM_11626_out0);
assign v$G1_8043_out0 = ((v$RD_6188_out0 && !v$RM_11628_out0) || (!v$RD_6188_out0) && v$RM_11628_out0);
assign v$G1_8045_out0 = ((v$RD_6190_out0 && !v$RM_11630_out0) || (!v$RD_6190_out0) && v$RM_11630_out0);
assign v$G1_8047_out0 = ((v$RD_6192_out0 && !v$RM_11632_out0) || (!v$RD_6192_out0) && v$RM_11632_out0);
assign v$G1_8049_out0 = ((v$RD_6194_out0 && !v$RM_11634_out0) || (!v$RD_6194_out0) && v$RM_11634_out0);
assign v$G1_8051_out0 = ((v$RD_6196_out0 && !v$RM_11636_out0) || (!v$RD_6196_out0) && v$RM_11636_out0);
assign v$G1_8053_out0 = ((v$RD_6198_out0 && !v$RM_11638_out0) || (!v$RD_6198_out0) && v$RM_11638_out0);
assign v$G1_8055_out0 = ((v$RD_6200_out0 && !v$RM_11640_out0) || (!v$RD_6200_out0) && v$RM_11640_out0);
assign v$G1_8490_out0 = ((v$RD_6635_out0 && !v$RM_12075_out0) || (!v$RD_6635_out0) && v$RM_12075_out0);
assign v$G1_8492_out0 = ((v$RD_6637_out0 && !v$RM_12077_out0) || (!v$RD_6637_out0) && v$RM_12077_out0);
assign v$G1_8496_out0 = ((v$RD_6641_out0 && !v$RM_12081_out0) || (!v$RD_6641_out0) && v$RM_12081_out0);
assign v$G1_8498_out0 = ((v$RD_6643_out0 && !v$RM_12083_out0) || (!v$RD_6643_out0) && v$RM_12083_out0);
assign v$G1_8500_out0 = ((v$RD_6645_out0 && !v$RM_12085_out0) || (!v$RD_6645_out0) && v$RM_12085_out0);
assign v$G1_8503_out0 = ((v$RD_6648_out0 && !v$RM_12088_out0) || (!v$RD_6648_out0) && v$RM_12088_out0);
assign v$G1_8505_out0 = ((v$RD_6650_out0 && !v$RM_12090_out0) || (!v$RD_6650_out0) && v$RM_12090_out0);
assign v$G1_8507_out0 = ((v$RD_6652_out0 && !v$RM_12092_out0) || (!v$RD_6652_out0) && v$RM_12092_out0);
assign v$G1_8509_out0 = ((v$RD_6654_out0 && !v$RM_12094_out0) || (!v$RD_6654_out0) && v$RM_12094_out0);
assign v$G1_8511_out0 = ((v$RD_6656_out0 && !v$RM_12096_out0) || (!v$RD_6656_out0) && v$RM_12096_out0);
assign v$G1_8513_out0 = ((v$RD_6658_out0 && !v$RM_12098_out0) || (!v$RD_6658_out0) && v$RM_12098_out0);
assign v$G1_8515_out0 = ((v$RD_6660_out0 && !v$RM_12100_out0) || (!v$RD_6660_out0) && v$RM_12100_out0);
assign v$G1_8517_out0 = ((v$RD_6662_out0 && !v$RM_12102_out0) || (!v$RD_6662_out0) && v$RM_12102_out0);
assign v$G1_8519_out0 = ((v$RD_6664_out0 && !v$RM_12104_out0) || (!v$RD_6664_out0) && v$RM_12104_out0);
assign v$S_9184_out0 = v$G1_8038_out0;
assign v$S_9648_out0 = v$G1_8502_out0;
assign v$G2_12562_out0 = v$RD_6171_out0 && v$RM_11611_out0;
assign v$G2_12564_out0 = v$RD_6173_out0 && v$RM_11613_out0;
assign v$G2_12568_out0 = v$RD_6177_out0 && v$RM_11617_out0;
assign v$G2_12570_out0 = v$RD_6179_out0 && v$RM_11619_out0;
assign v$G2_12572_out0 = v$RD_6181_out0 && v$RM_11621_out0;
assign v$G2_12575_out0 = v$RD_6184_out0 && v$RM_11624_out0;
assign v$G2_12577_out0 = v$RD_6186_out0 && v$RM_11626_out0;
assign v$G2_12579_out0 = v$RD_6188_out0 && v$RM_11628_out0;
assign v$G2_12581_out0 = v$RD_6190_out0 && v$RM_11630_out0;
assign v$G2_12583_out0 = v$RD_6192_out0 && v$RM_11632_out0;
assign v$G2_12585_out0 = v$RD_6194_out0 && v$RM_11634_out0;
assign v$G2_12587_out0 = v$RD_6196_out0 && v$RM_11636_out0;
assign v$G2_12589_out0 = v$RD_6198_out0 && v$RM_11638_out0;
assign v$G2_12591_out0 = v$RD_6200_out0 && v$RM_11640_out0;
assign v$G2_13026_out0 = v$RD_6635_out0 && v$RM_12075_out0;
assign v$G2_13028_out0 = v$RD_6637_out0 && v$RM_12077_out0;
assign v$G2_13032_out0 = v$RD_6641_out0 && v$RM_12081_out0;
assign v$G2_13034_out0 = v$RD_6643_out0 && v$RM_12083_out0;
assign v$G2_13036_out0 = v$RD_6645_out0 && v$RM_12085_out0;
assign v$G2_13039_out0 = v$RD_6648_out0 && v$RM_12088_out0;
assign v$G2_13041_out0 = v$RD_6650_out0 && v$RM_12090_out0;
assign v$G2_13043_out0 = v$RD_6652_out0 && v$RM_12092_out0;
assign v$G2_13045_out0 = v$RD_6654_out0 && v$RM_12094_out0;
assign v$G2_13047_out0 = v$RD_6656_out0 && v$RM_12096_out0;
assign v$G2_13049_out0 = v$RD_6658_out0 && v$RM_12098_out0;
assign v$G2_13051_out0 = v$RD_6660_out0 && v$RM_12100_out0;
assign v$G2_13053_out0 = v$RD_6662_out0 && v$RM_12102_out0;
assign v$G2_13055_out0 = v$RD_6664_out0 && v$RM_12104_out0;
assign v$S_4675_out0 = v$S_9184_out0;
assign v$S_4690_out0 = v$S_9648_out0;
assign v$CARRY_5171_out0 = v$G2_12562_out0;
assign v$CARRY_5173_out0 = v$G2_12564_out0;
assign v$CARRY_5177_out0 = v$G2_12568_out0;
assign v$CARRY_5179_out0 = v$G2_12570_out0;
assign v$CARRY_5181_out0 = v$G2_12572_out0;
assign v$CARRY_5184_out0 = v$G2_12575_out0;
assign v$CARRY_5186_out0 = v$G2_12577_out0;
assign v$CARRY_5188_out0 = v$G2_12579_out0;
assign v$CARRY_5190_out0 = v$G2_12581_out0;
assign v$CARRY_5192_out0 = v$G2_12583_out0;
assign v$CARRY_5194_out0 = v$G2_12585_out0;
assign v$CARRY_5196_out0 = v$G2_12587_out0;
assign v$CARRY_5198_out0 = v$G2_12589_out0;
assign v$CARRY_5200_out0 = v$G2_12591_out0;
assign v$CARRY_5635_out0 = v$G2_13026_out0;
assign v$CARRY_5637_out0 = v$G2_13028_out0;
assign v$CARRY_5641_out0 = v$G2_13032_out0;
assign v$CARRY_5643_out0 = v$G2_13034_out0;
assign v$CARRY_5645_out0 = v$G2_13036_out0;
assign v$CARRY_5648_out0 = v$G2_13039_out0;
assign v$CARRY_5650_out0 = v$G2_13041_out0;
assign v$CARRY_5652_out0 = v$G2_13043_out0;
assign v$CARRY_5654_out0 = v$G2_13045_out0;
assign v$CARRY_5656_out0 = v$G2_13047_out0;
assign v$CARRY_5658_out0 = v$G2_13049_out0;
assign v$CARRY_5660_out0 = v$G2_13051_out0;
assign v$CARRY_5662_out0 = v$G2_13053_out0;
assign v$CARRY_5664_out0 = v$G2_13055_out0;
assign v$S_9172_out0 = v$G1_8026_out0;
assign v$S_9174_out0 = v$G1_8028_out0;
assign v$S_9178_out0 = v$G1_8032_out0;
assign v$S_9180_out0 = v$G1_8034_out0;
assign v$S_9182_out0 = v$G1_8036_out0;
assign v$S_9185_out0 = v$G1_8039_out0;
assign v$S_9187_out0 = v$G1_8041_out0;
assign v$S_9189_out0 = v$G1_8043_out0;
assign v$S_9191_out0 = v$G1_8045_out0;
assign v$S_9193_out0 = v$G1_8047_out0;
assign v$S_9195_out0 = v$G1_8049_out0;
assign v$S_9197_out0 = v$G1_8051_out0;
assign v$S_9199_out0 = v$G1_8053_out0;
assign v$S_9201_out0 = v$G1_8055_out0;
assign v$S_9636_out0 = v$G1_8490_out0;
assign v$S_9638_out0 = v$G1_8492_out0;
assign v$S_9642_out0 = v$G1_8496_out0;
assign v$S_9644_out0 = v$G1_8498_out0;
assign v$S_9646_out0 = v$G1_8500_out0;
assign v$S_9649_out0 = v$G1_8503_out0;
assign v$S_9651_out0 = v$G1_8505_out0;
assign v$S_9653_out0 = v$G1_8507_out0;
assign v$S_9655_out0 = v$G1_8509_out0;
assign v$S_9657_out0 = v$G1_8511_out0;
assign v$S_9659_out0 = v$G1_8513_out0;
assign v$S_9661_out0 = v$G1_8515_out0;
assign v$S_9663_out0 = v$G1_8517_out0;
assign v$S_9665_out0 = v$G1_8519_out0;
assign v$CIN_9965_out0 = v$CARRY_5183_out0;
assign v$CIN_10189_out0 = v$CARRY_5647_out0;
assign v$_56_out0 = { v$_2392_out0,v$S_4675_out0 };
assign v$_57_out0 = { v$_2393_out0,v$S_4690_out0 };
assign v$RD_6189_out0 = v$CIN_9965_out0;
assign v$RD_6653_out0 = v$CIN_10189_out0;
assign v$RM_11612_out0 = v$S_9172_out0;
assign v$RM_11614_out0 = v$S_9174_out0;
assign v$RM_11618_out0 = v$S_9178_out0;
assign v$RM_11620_out0 = v$S_9180_out0;
assign v$RM_11622_out0 = v$S_9182_out0;
assign v$RM_11625_out0 = v$S_9185_out0;
assign v$RM_11627_out0 = v$S_9187_out0;
assign v$RM_11629_out0 = v$S_9189_out0;
assign v$RM_11631_out0 = v$S_9191_out0;
assign v$RM_11633_out0 = v$S_9193_out0;
assign v$RM_11635_out0 = v$S_9195_out0;
assign v$RM_11637_out0 = v$S_9197_out0;
assign v$RM_11639_out0 = v$S_9199_out0;
assign v$RM_11641_out0 = v$S_9201_out0;
assign v$RM_12076_out0 = v$S_9636_out0;
assign v$RM_12078_out0 = v$S_9638_out0;
assign v$RM_12082_out0 = v$S_9642_out0;
assign v$RM_12084_out0 = v$S_9644_out0;
assign v$RM_12086_out0 = v$S_9646_out0;
assign v$RM_12089_out0 = v$S_9649_out0;
assign v$RM_12091_out0 = v$S_9651_out0;
assign v$RM_12093_out0 = v$S_9653_out0;
assign v$RM_12095_out0 = v$S_9655_out0;
assign v$RM_12097_out0 = v$S_9657_out0;
assign v$RM_12099_out0 = v$S_9659_out0;
assign v$RM_12101_out0 = v$S_9661_out0;
assign v$RM_12103_out0 = v$S_9663_out0;
assign v$RM_12105_out0 = v$S_9665_out0;
assign v$G1_8044_out0 = ((v$RD_6189_out0 && !v$RM_11629_out0) || (!v$RD_6189_out0) && v$RM_11629_out0);
assign v$G1_8508_out0 = ((v$RD_6653_out0 && !v$RM_12093_out0) || (!v$RD_6653_out0) && v$RM_12093_out0);
assign v$G2_12580_out0 = v$RD_6189_out0 && v$RM_11629_out0;
assign v$G2_13044_out0 = v$RD_6653_out0 && v$RM_12093_out0;
assign v$CARRY_5189_out0 = v$G2_12580_out0;
assign v$CARRY_5653_out0 = v$G2_13044_out0;
assign v$S_9190_out0 = v$G1_8044_out0;
assign v$S_9654_out0 = v$G1_8508_out0;
assign v$S_1376_out0 = v$S_9190_out0;
assign v$S_1600_out0 = v$S_9654_out0;
assign v$G1_4152_out0 = v$CARRY_5189_out0 || v$CARRY_5188_out0;
assign v$G1_4376_out0 = v$CARRY_5653_out0 || v$CARRY_5652_out0;
assign v$COUT_844_out0 = v$G1_4152_out0;
assign v$COUT_1068_out0 = v$G1_4376_out0;
assign v$CIN_9971_out0 = v$COUT_844_out0;
assign v$CIN_10195_out0 = v$COUT_1068_out0;
assign v$RD_6201_out0 = v$CIN_9971_out0;
assign v$RD_6665_out0 = v$CIN_10195_out0;
assign v$G1_8056_out0 = ((v$RD_6201_out0 && !v$RM_11641_out0) || (!v$RD_6201_out0) && v$RM_11641_out0);
assign v$G1_8520_out0 = ((v$RD_6665_out0 && !v$RM_12105_out0) || (!v$RD_6665_out0) && v$RM_12105_out0);
assign v$G2_12592_out0 = v$RD_6201_out0 && v$RM_11641_out0;
assign v$G2_13056_out0 = v$RD_6665_out0 && v$RM_12105_out0;
assign v$CARRY_5201_out0 = v$G2_12592_out0;
assign v$CARRY_5665_out0 = v$G2_13056_out0;
assign v$S_9202_out0 = v$G1_8056_out0;
assign v$S_9666_out0 = v$G1_8520_out0;
assign v$S_1382_out0 = v$S_9202_out0;
assign v$S_1606_out0 = v$S_9666_out0;
assign v$G1_4158_out0 = v$CARRY_5201_out0 || v$CARRY_5200_out0;
assign v$G1_4382_out0 = v$CARRY_5665_out0 || v$CARRY_5664_out0;
assign v$COUT_850_out0 = v$G1_4158_out0;
assign v$COUT_1074_out0 = v$G1_4382_out0;
assign v$_4792_out0 = { v$S_1376_out0,v$S_1382_out0 };
assign v$_4807_out0 = { v$S_1600_out0,v$S_1606_out0 };
assign v$CIN_9966_out0 = v$COUT_850_out0;
assign v$CIN_10190_out0 = v$COUT_1074_out0;
assign v$RD_6191_out0 = v$CIN_9966_out0;
assign v$RD_6655_out0 = v$CIN_10190_out0;
assign v$G1_8046_out0 = ((v$RD_6191_out0 && !v$RM_11631_out0) || (!v$RD_6191_out0) && v$RM_11631_out0);
assign v$G1_8510_out0 = ((v$RD_6655_out0 && !v$RM_12095_out0) || (!v$RD_6655_out0) && v$RM_12095_out0);
assign v$G2_12582_out0 = v$RD_6191_out0 && v$RM_11631_out0;
assign v$G2_13046_out0 = v$RD_6655_out0 && v$RM_12095_out0;
assign v$CARRY_5191_out0 = v$G2_12582_out0;
assign v$CARRY_5655_out0 = v$G2_13046_out0;
assign v$S_9192_out0 = v$G1_8046_out0;
assign v$S_9656_out0 = v$G1_8510_out0;
assign v$S_1377_out0 = v$S_9192_out0;
assign v$S_1601_out0 = v$S_9656_out0;
assign v$G1_4153_out0 = v$CARRY_5191_out0 || v$CARRY_5190_out0;
assign v$G1_4377_out0 = v$CARRY_5655_out0 || v$CARRY_5654_out0;
assign v$COUT_845_out0 = v$G1_4153_out0;
assign v$COUT_1069_out0 = v$G1_4377_out0;
assign v$_2562_out0 = { v$_4792_out0,v$S_1377_out0 };
assign v$_2577_out0 = { v$_4807_out0,v$S_1601_out0 };
assign v$CIN_9961_out0 = v$COUT_845_out0;
assign v$CIN_10185_out0 = v$COUT_1069_out0;
assign v$RD_6180_out0 = v$CIN_9961_out0;
assign v$RD_6644_out0 = v$CIN_10185_out0;
assign v$G1_8035_out0 = ((v$RD_6180_out0 && !v$RM_11620_out0) || (!v$RD_6180_out0) && v$RM_11620_out0);
assign v$G1_8499_out0 = ((v$RD_6644_out0 && !v$RM_12084_out0) || (!v$RD_6644_out0) && v$RM_12084_out0);
assign v$G2_12571_out0 = v$RD_6180_out0 && v$RM_11620_out0;
assign v$G2_13035_out0 = v$RD_6644_out0 && v$RM_12084_out0;
assign v$CARRY_5180_out0 = v$G2_12571_out0;
assign v$CARRY_5644_out0 = v$G2_13035_out0;
assign v$S_9181_out0 = v$G1_8035_out0;
assign v$S_9645_out0 = v$G1_8499_out0;
assign v$S_1372_out0 = v$S_9181_out0;
assign v$S_1596_out0 = v$S_9645_out0;
assign v$G1_4148_out0 = v$CARRY_5180_out0 || v$CARRY_5179_out0;
assign v$G1_4372_out0 = v$CARRY_5644_out0 || v$CARRY_5643_out0;
assign v$COUT_840_out0 = v$G1_4148_out0;
assign v$COUT_1064_out0 = v$G1_4372_out0;
assign v$_7042_out0 = { v$_2562_out0,v$S_1372_out0 };
assign v$_7057_out0 = { v$_2577_out0,v$S_1596_out0 };
assign v$CIN_9960_out0 = v$COUT_840_out0;
assign v$CIN_10184_out0 = v$COUT_1064_out0;
assign v$RD_6178_out0 = v$CIN_9960_out0;
assign v$RD_6642_out0 = v$CIN_10184_out0;
assign v$G1_8033_out0 = ((v$RD_6178_out0 && !v$RM_11618_out0) || (!v$RD_6178_out0) && v$RM_11618_out0);
assign v$G1_8497_out0 = ((v$RD_6642_out0 && !v$RM_12082_out0) || (!v$RD_6642_out0) && v$RM_12082_out0);
assign v$G2_12569_out0 = v$RD_6178_out0 && v$RM_11618_out0;
assign v$G2_13033_out0 = v$RD_6642_out0 && v$RM_12082_out0;
assign v$CARRY_5178_out0 = v$G2_12569_out0;
assign v$CARRY_5642_out0 = v$G2_13033_out0;
assign v$S_9179_out0 = v$G1_8033_out0;
assign v$S_9643_out0 = v$G1_8497_out0;
assign v$S_1371_out0 = v$S_9179_out0;
assign v$S_1595_out0 = v$S_9643_out0;
assign v$G1_4147_out0 = v$CARRY_5178_out0 || v$CARRY_5177_out0;
assign v$G1_4371_out0 = v$CARRY_5642_out0 || v$CARRY_5641_out0;
assign v$COUT_839_out0 = v$G1_4147_out0;
assign v$COUT_1063_out0 = v$G1_4371_out0;
assign v$_13528_out0 = { v$_7042_out0,v$S_1371_out0 };
assign v$_13543_out0 = { v$_7057_out0,v$S_1595_out0 };
assign v$CIN_9967_out0 = v$COUT_839_out0;
assign v$CIN_10191_out0 = v$COUT_1063_out0;
assign v$RD_6193_out0 = v$CIN_9967_out0;
assign v$RD_6657_out0 = v$CIN_10191_out0;
assign v$G1_8048_out0 = ((v$RD_6193_out0 && !v$RM_11633_out0) || (!v$RD_6193_out0) && v$RM_11633_out0);
assign v$G1_8512_out0 = ((v$RD_6657_out0 && !v$RM_12097_out0) || (!v$RD_6657_out0) && v$RM_12097_out0);
assign v$G2_12584_out0 = v$RD_6193_out0 && v$RM_11633_out0;
assign v$G2_13048_out0 = v$RD_6657_out0 && v$RM_12097_out0;
assign v$CARRY_5193_out0 = v$G2_12584_out0;
assign v$CARRY_5657_out0 = v$G2_13048_out0;
assign v$S_9194_out0 = v$G1_8048_out0;
assign v$S_9658_out0 = v$G1_8512_out0;
assign v$S_1378_out0 = v$S_9194_out0;
assign v$S_1602_out0 = v$S_9658_out0;
assign v$G1_4154_out0 = v$CARRY_5193_out0 || v$CARRY_5192_out0;
assign v$G1_4378_out0 = v$CARRY_5657_out0 || v$CARRY_5656_out0;
assign v$COUT_846_out0 = v$G1_4154_out0;
assign v$COUT_1070_out0 = v$G1_4378_out0;
assign v$_3321_out0 = { v$_13528_out0,v$S_1378_out0 };
assign v$_3336_out0 = { v$_13543_out0,v$S_1602_out0 };
assign v$CIN_9968_out0 = v$COUT_846_out0;
assign v$CIN_10192_out0 = v$COUT_1070_out0;
assign v$RD_6195_out0 = v$CIN_9968_out0;
assign v$RD_6659_out0 = v$CIN_10192_out0;
assign v$G1_8050_out0 = ((v$RD_6195_out0 && !v$RM_11635_out0) || (!v$RD_6195_out0) && v$RM_11635_out0);
assign v$G1_8514_out0 = ((v$RD_6659_out0 && !v$RM_12099_out0) || (!v$RD_6659_out0) && v$RM_12099_out0);
assign v$G2_12586_out0 = v$RD_6195_out0 && v$RM_11635_out0;
assign v$G2_13050_out0 = v$RD_6659_out0 && v$RM_12099_out0;
assign v$CARRY_5195_out0 = v$G2_12586_out0;
assign v$CARRY_5659_out0 = v$G2_13050_out0;
assign v$S_9196_out0 = v$G1_8050_out0;
assign v$S_9660_out0 = v$G1_8514_out0;
assign v$S_1379_out0 = v$S_9196_out0;
assign v$S_1603_out0 = v$S_9660_out0;
assign v$G1_4155_out0 = v$CARRY_5195_out0 || v$CARRY_5194_out0;
assign v$G1_4379_out0 = v$CARRY_5659_out0 || v$CARRY_5658_out0;
assign v$COUT_847_out0 = v$G1_4155_out0;
assign v$COUT_1071_out0 = v$G1_4379_out0;
assign v$_7157_out0 = { v$_3321_out0,v$S_1379_out0 };
assign v$_7172_out0 = { v$_3336_out0,v$S_1603_out0 };
assign v$CIN_9970_out0 = v$COUT_847_out0;
assign v$CIN_10194_out0 = v$COUT_1071_out0;
assign v$RD_6199_out0 = v$CIN_9970_out0;
assign v$RD_6663_out0 = v$CIN_10194_out0;
assign v$G1_8054_out0 = ((v$RD_6199_out0 && !v$RM_11639_out0) || (!v$RD_6199_out0) && v$RM_11639_out0);
assign v$G1_8518_out0 = ((v$RD_6663_out0 && !v$RM_12103_out0) || (!v$RD_6663_out0) && v$RM_12103_out0);
assign v$G2_12590_out0 = v$RD_6199_out0 && v$RM_11639_out0;
assign v$G2_13054_out0 = v$RD_6663_out0 && v$RM_12103_out0;
assign v$CARRY_5199_out0 = v$G2_12590_out0;
assign v$CARRY_5663_out0 = v$G2_13054_out0;
assign v$S_9200_out0 = v$G1_8054_out0;
assign v$S_9664_out0 = v$G1_8518_out0;
assign v$S_1381_out0 = v$S_9200_out0;
assign v$S_1605_out0 = v$S_9664_out0;
assign v$G1_4157_out0 = v$CARRY_5199_out0 || v$CARRY_5198_out0;
assign v$G1_4381_out0 = v$CARRY_5663_out0 || v$CARRY_5662_out0;
assign v$COUT_849_out0 = v$G1_4157_out0;
assign v$COUT_1073_out0 = v$G1_4381_out0;
assign v$_4759_out0 = { v$_7157_out0,v$S_1381_out0 };
assign v$_4774_out0 = { v$_7172_out0,v$S_1605_out0 };
assign v$CIN_9963_out0 = v$COUT_849_out0;
assign v$CIN_10187_out0 = v$COUT_1073_out0;
assign v$RD_6185_out0 = v$CIN_9963_out0;
assign v$RD_6649_out0 = v$CIN_10187_out0;
assign v$G1_8040_out0 = ((v$RD_6185_out0 && !v$RM_11625_out0) || (!v$RD_6185_out0) && v$RM_11625_out0);
assign v$G1_8504_out0 = ((v$RD_6649_out0 && !v$RM_12089_out0) || (!v$RD_6649_out0) && v$RM_12089_out0);
assign v$G2_12576_out0 = v$RD_6185_out0 && v$RM_11625_out0;
assign v$G2_13040_out0 = v$RD_6649_out0 && v$RM_12089_out0;
assign v$CARRY_5185_out0 = v$G2_12576_out0;
assign v$CARRY_5649_out0 = v$G2_13040_out0;
assign v$S_9186_out0 = v$G1_8040_out0;
assign v$S_9650_out0 = v$G1_8504_out0;
assign v$S_1374_out0 = v$S_9186_out0;
assign v$S_1598_out0 = v$S_9650_out0;
assign v$G1_4150_out0 = v$CARRY_5185_out0 || v$CARRY_5184_out0;
assign v$G1_4374_out0 = v$CARRY_5649_out0 || v$CARRY_5648_out0;
assign v$COUT_842_out0 = v$G1_4150_out0;
assign v$COUT_1066_out0 = v$G1_4374_out0;
assign v$_6936_out0 = { v$_4759_out0,v$S_1374_out0 };
assign v$_6951_out0 = { v$_4774_out0,v$S_1598_out0 };
assign v$CIN_9964_out0 = v$COUT_842_out0;
assign v$CIN_10188_out0 = v$COUT_1066_out0;
assign v$RD_6187_out0 = v$CIN_9964_out0;
assign v$RD_6651_out0 = v$CIN_10188_out0;
assign v$G1_8042_out0 = ((v$RD_6187_out0 && !v$RM_11627_out0) || (!v$RD_6187_out0) && v$RM_11627_out0);
assign v$G1_8506_out0 = ((v$RD_6651_out0 && !v$RM_12091_out0) || (!v$RD_6651_out0) && v$RM_12091_out0);
assign v$G2_12578_out0 = v$RD_6187_out0 && v$RM_11627_out0;
assign v$G2_13042_out0 = v$RD_6651_out0 && v$RM_12091_out0;
assign v$CARRY_5187_out0 = v$G2_12578_out0;
assign v$CARRY_5651_out0 = v$G2_13042_out0;
assign v$S_9188_out0 = v$G1_8042_out0;
assign v$S_9652_out0 = v$G1_8506_out0;
assign v$S_1375_out0 = v$S_9188_out0;
assign v$S_1599_out0 = v$S_9652_out0;
assign v$G1_4151_out0 = v$CARRY_5187_out0 || v$CARRY_5186_out0;
assign v$G1_4375_out0 = v$CARRY_5651_out0 || v$CARRY_5650_out0;
assign v$COUT_843_out0 = v$G1_4151_out0;
assign v$COUT_1067_out0 = v$G1_4375_out0;
assign v$_5812_out0 = { v$_6936_out0,v$S_1375_out0 };
assign v$_5827_out0 = { v$_6951_out0,v$S_1599_out0 };
assign v$CIN_9969_out0 = v$COUT_843_out0;
assign v$CIN_10193_out0 = v$COUT_1067_out0;
assign v$RD_6197_out0 = v$CIN_9969_out0;
assign v$RD_6661_out0 = v$CIN_10193_out0;
assign v$G1_8052_out0 = ((v$RD_6197_out0 && !v$RM_11637_out0) || (!v$RD_6197_out0) && v$RM_11637_out0);
assign v$G1_8516_out0 = ((v$RD_6661_out0 && !v$RM_12101_out0) || (!v$RD_6661_out0) && v$RM_12101_out0);
assign v$G2_12588_out0 = v$RD_6197_out0 && v$RM_11637_out0;
assign v$G2_13052_out0 = v$RD_6661_out0 && v$RM_12101_out0;
assign v$CARRY_5197_out0 = v$G2_12588_out0;
assign v$CARRY_5661_out0 = v$G2_13052_out0;
assign v$S_9198_out0 = v$G1_8052_out0;
assign v$S_9662_out0 = v$G1_8516_out0;
assign v$S_1380_out0 = v$S_9198_out0;
assign v$S_1604_out0 = v$S_9662_out0;
assign v$G1_4156_out0 = v$CARRY_5197_out0 || v$CARRY_5196_out0;
assign v$G1_4380_out0 = v$CARRY_5661_out0 || v$CARRY_5660_out0;
assign v$COUT_848_out0 = v$G1_4156_out0;
assign v$COUT_1072_out0 = v$G1_4380_out0;
assign v$_2036_out0 = { v$_5812_out0,v$S_1380_out0 };
assign v$_2051_out0 = { v$_5827_out0,v$S_1604_out0 };
assign v$CIN_9957_out0 = v$COUT_848_out0;
assign v$CIN_10181_out0 = v$COUT_1072_out0;
assign v$RD_6172_out0 = v$CIN_9957_out0;
assign v$RD_6636_out0 = v$CIN_10181_out0;
assign v$G1_8027_out0 = ((v$RD_6172_out0 && !v$RM_11612_out0) || (!v$RD_6172_out0) && v$RM_11612_out0);
assign v$G1_8491_out0 = ((v$RD_6636_out0 && !v$RM_12076_out0) || (!v$RD_6636_out0) && v$RM_12076_out0);
assign v$G2_12563_out0 = v$RD_6172_out0 && v$RM_11612_out0;
assign v$G2_13027_out0 = v$RD_6636_out0 && v$RM_12076_out0;
assign v$CARRY_5172_out0 = v$G2_12563_out0;
assign v$CARRY_5636_out0 = v$G2_13027_out0;
assign v$S_9173_out0 = v$G1_8027_out0;
assign v$S_9637_out0 = v$G1_8491_out0;
assign v$S_1368_out0 = v$S_9173_out0;
assign v$S_1592_out0 = v$S_9637_out0;
assign v$G1_4144_out0 = v$CARRY_5172_out0 || v$CARRY_5171_out0;
assign v$G1_4368_out0 = v$CARRY_5636_out0 || v$CARRY_5635_out0;
assign v$COUT_836_out0 = v$G1_4144_out0;
assign v$COUT_1060_out0 = v$G1_4368_out0;
assign v$_2803_out0 = { v$_2036_out0,v$S_1368_out0 };
assign v$_2818_out0 = { v$_2051_out0,v$S_1592_out0 };
assign v$CIN_9962_out0 = v$COUT_836_out0;
assign v$CIN_10186_out0 = v$COUT_1060_out0;
assign v$RD_6182_out0 = v$CIN_9962_out0;
assign v$RD_6646_out0 = v$CIN_10186_out0;
assign v$G1_8037_out0 = ((v$RD_6182_out0 && !v$RM_11622_out0) || (!v$RD_6182_out0) && v$RM_11622_out0);
assign v$G1_8501_out0 = ((v$RD_6646_out0 && !v$RM_12086_out0) || (!v$RD_6646_out0) && v$RM_12086_out0);
assign v$G2_12573_out0 = v$RD_6182_out0 && v$RM_11622_out0;
assign v$G2_13037_out0 = v$RD_6646_out0 && v$RM_12086_out0;
assign v$CARRY_5182_out0 = v$G2_12573_out0;
assign v$CARRY_5646_out0 = v$G2_13037_out0;
assign v$S_9183_out0 = v$G1_8037_out0;
assign v$S_9647_out0 = v$G1_8501_out0;
assign v$S_1373_out0 = v$S_9183_out0;
assign v$S_1597_out0 = v$S_9647_out0;
assign v$G1_4149_out0 = v$CARRY_5182_out0 || v$CARRY_5181_out0;
assign v$G1_4373_out0 = v$CARRY_5646_out0 || v$CARRY_5645_out0;
assign v$COUT_841_out0 = v$G1_4149_out0;
assign v$COUT_1065_out0 = v$G1_4373_out0;
assign v$_1835_out0 = { v$_2803_out0,v$S_1373_out0 };
assign v$_1850_out0 = { v$_2818_out0,v$S_1597_out0 };
assign v$CIN_9958_out0 = v$COUT_841_out0;
assign v$CIN_10182_out0 = v$COUT_1065_out0;
assign v$RD_6174_out0 = v$CIN_9958_out0;
assign v$RD_6638_out0 = v$CIN_10182_out0;
assign v$G1_8029_out0 = ((v$RD_6174_out0 && !v$RM_11614_out0) || (!v$RD_6174_out0) && v$RM_11614_out0);
assign v$G1_8493_out0 = ((v$RD_6638_out0 && !v$RM_12078_out0) || (!v$RD_6638_out0) && v$RM_12078_out0);
assign v$G2_12565_out0 = v$RD_6174_out0 && v$RM_11614_out0;
assign v$G2_13029_out0 = v$RD_6638_out0 && v$RM_12078_out0;
assign v$CARRY_5174_out0 = v$G2_12565_out0;
assign v$CARRY_5638_out0 = v$G2_13029_out0;
assign v$S_9175_out0 = v$G1_8029_out0;
assign v$S_9639_out0 = v$G1_8493_out0;
assign v$S_1369_out0 = v$S_9175_out0;
assign v$S_1593_out0 = v$S_9639_out0;
assign v$G1_4145_out0 = v$CARRY_5174_out0 || v$CARRY_5173_out0;
assign v$G1_4369_out0 = v$CARRY_5638_out0 || v$CARRY_5637_out0;
assign v$COUT_837_out0 = v$G1_4145_out0;
assign v$COUT_1061_out0 = v$G1_4369_out0;
assign v$_4559_out0 = { v$_1835_out0,v$S_1369_out0 };
assign v$_4574_out0 = { v$_1850_out0,v$S_1593_out0 };
assign v$RM_3506_out0 = v$COUT_837_out0;
assign v$RM_3730_out0 = v$COUT_1061_out0;
assign v$RM_11615_out0 = v$RM_3506_out0;
assign v$RM_12079_out0 = v$RM_3730_out0;
assign v$G1_8030_out0 = ((v$RD_6175_out0 && !v$RM_11615_out0) || (!v$RD_6175_out0) && v$RM_11615_out0);
assign v$G1_8494_out0 = ((v$RD_6639_out0 && !v$RM_12079_out0) || (!v$RD_6639_out0) && v$RM_12079_out0);
assign v$G2_12566_out0 = v$RD_6175_out0 && v$RM_11615_out0;
assign v$G2_13030_out0 = v$RD_6639_out0 && v$RM_12079_out0;
assign v$CARRY_5175_out0 = v$G2_12566_out0;
assign v$CARRY_5639_out0 = v$G2_13030_out0;
assign v$S_9176_out0 = v$G1_8030_out0;
assign v$S_9640_out0 = v$G1_8494_out0;
assign v$RM_11616_out0 = v$S_9176_out0;
assign v$RM_12080_out0 = v$S_9640_out0;
assign v$G1_8031_out0 = ((v$RD_6176_out0 && !v$RM_11616_out0) || (!v$RD_6176_out0) && v$RM_11616_out0);
assign v$G1_8495_out0 = ((v$RD_6640_out0 && !v$RM_12080_out0) || (!v$RD_6640_out0) && v$RM_12080_out0);
assign v$G2_12567_out0 = v$RD_6176_out0 && v$RM_11616_out0;
assign v$G2_13031_out0 = v$RD_6640_out0 && v$RM_12080_out0;
assign v$CARRY_5176_out0 = v$G2_12567_out0;
assign v$CARRY_5640_out0 = v$G2_13031_out0;
assign v$S_9177_out0 = v$G1_8031_out0;
assign v$S_9641_out0 = v$G1_8495_out0;
assign v$S_1370_out0 = v$S_9177_out0;
assign v$S_1594_out0 = v$S_9641_out0;
assign v$G1_4146_out0 = v$CARRY_5176_out0 || v$CARRY_5175_out0;
assign v$G1_4370_out0 = v$CARRY_5640_out0 || v$CARRY_5639_out0;
assign v$COUT_838_out0 = v$G1_4146_out0;
assign v$COUT_1062_out0 = v$G1_4370_out0;
assign v$_10661_out0 = { v$_4559_out0,v$S_1370_out0 };
assign v$_10676_out0 = { v$_4574_out0,v$S_1594_out0 };
assign v$_10956_out0 = { v$_10661_out0,v$COUT_838_out0 };
assign v$_10971_out0 = { v$_10676_out0,v$COUT_1062_out0 };
assign v$COUT_10926_out0 = v$_10956_out0;
assign v$COUT_10941_out0 = v$_10971_out0;
assign v$CIN_2368_out0 = v$COUT_10926_out0;
assign v$CIN_2383_out0 = v$COUT_10941_out0;
assign v$_481_out0 = v$CIN_2368_out0[8:8];
assign v$_496_out0 = v$CIN_2383_out0[8:8];
assign v$_1786_out0 = v$CIN_2368_out0[6:6];
assign v$_1801_out0 = v$CIN_2383_out0[6:6];
assign v$_2168_out0 = v$CIN_2368_out0[3:3];
assign v$_2183_out0 = v$CIN_2383_out0[3:3];
assign v$_2207_out0 = v$CIN_2368_out0[15:15];
assign v$_2221_out0 = v$CIN_2383_out0[15:15];
assign v$_2515_out0 = v$CIN_2368_out0[0:0];
assign v$_2530_out0 = v$CIN_2383_out0[0:0];
assign v$_3064_out0 = v$CIN_2368_out0[9:9];
assign v$_3079_out0 = v$CIN_2383_out0[9:9];
assign v$_3098_out0 = v$CIN_2368_out0[2:2];
assign v$_3113_out0 = v$CIN_2383_out0[2:2];
assign v$_3152_out0 = v$CIN_2368_out0[7:7];
assign v$_3167_out0 = v$CIN_2383_out0[7:7];
assign v$_3836_out0 = v$CIN_2368_out0[1:1];
assign v$_3851_out0 = v$CIN_2383_out0[1:1];
assign v$_3874_out0 = v$CIN_2368_out0[10:10];
assign v$_3889_out0 = v$CIN_2383_out0[10:10];
assign v$_6813_out0 = v$CIN_2368_out0[11:11];
assign v$_6828_out0 = v$CIN_2383_out0[11:11];
assign v$_7657_out0 = v$CIN_2368_out0[12:12];
assign v$_7672_out0 = v$CIN_2383_out0[12:12];
assign v$_8712_out0 = v$CIN_2368_out0[13:13];
assign v$_8727_out0 = v$CIN_2383_out0[13:13];
assign v$_8782_out0 = v$CIN_2368_out0[14:14];
assign v$_8797_out0 = v$CIN_2383_out0[14:14];
assign v$_10732_out0 = v$CIN_2368_out0[5:5];
assign v$_10747_out0 = v$CIN_2383_out0[5:5];
assign v$_13461_out0 = v$CIN_2368_out0[4:4];
assign v$_13476_out0 = v$CIN_2383_out0[4:4];
assign v$RM_3549_out0 = v$_7657_out0;
assign v$RM_3550_out0 = v$_8782_out0;
assign v$RM_3552_out0 = v$_10732_out0;
assign v$RM_3553_out0 = v$_13461_out0;
assign v$RM_3554_out0 = v$_8712_out0;
assign v$RM_3555_out0 = v$_3064_out0;
assign v$RM_3556_out0 = v$_3874_out0;
assign v$RM_3557_out0 = v$_3836_out0;
assign v$RM_3558_out0 = v$_2168_out0;
assign v$RM_3559_out0 = v$_1786_out0;
assign v$RM_3560_out0 = v$_3152_out0;
assign v$RM_3561_out0 = v$_6813_out0;
assign v$RM_3562_out0 = v$_481_out0;
assign v$RM_3563_out0 = v$_3098_out0;
assign v$RM_3773_out0 = v$_7672_out0;
assign v$RM_3774_out0 = v$_8797_out0;
assign v$RM_3776_out0 = v$_10747_out0;
assign v$RM_3777_out0 = v$_13476_out0;
assign v$RM_3778_out0 = v$_8727_out0;
assign v$RM_3779_out0 = v$_3079_out0;
assign v$RM_3780_out0 = v$_3889_out0;
assign v$RM_3781_out0 = v$_3851_out0;
assign v$RM_3782_out0 = v$_2183_out0;
assign v$RM_3783_out0 = v$_1801_out0;
assign v$RM_3784_out0 = v$_3167_out0;
assign v$RM_3785_out0 = v$_6828_out0;
assign v$RM_3786_out0 = v$_496_out0;
assign v$RM_3787_out0 = v$_3113_out0;
assign v$CIN_10004_out0 = v$_2207_out0;
assign v$CIN_10228_out0 = v$_2221_out0;
assign v$RM_11716_out0 = v$_2515_out0;
assign v$RM_12180_out0 = v$_2530_out0;
assign v$RD_6269_out0 = v$CIN_10004_out0;
assign v$RD_6733_out0 = v$CIN_10228_out0;
assign v$G1_8131_out0 = ((v$RD_6276_out0 && !v$RM_11716_out0) || (!v$RD_6276_out0) && v$RM_11716_out0);
assign v$G1_8595_out0 = ((v$RD_6740_out0 && !v$RM_12180_out0) || (!v$RD_6740_out0) && v$RM_12180_out0);
assign v$RM_11704_out0 = v$RM_3549_out0;
assign v$RM_11706_out0 = v$RM_3550_out0;
assign v$RM_11710_out0 = v$RM_3552_out0;
assign v$RM_11712_out0 = v$RM_3553_out0;
assign v$RM_11714_out0 = v$RM_3554_out0;
assign v$RM_11717_out0 = v$RM_3555_out0;
assign v$RM_11719_out0 = v$RM_3556_out0;
assign v$RM_11721_out0 = v$RM_3557_out0;
assign v$RM_11723_out0 = v$RM_3558_out0;
assign v$RM_11725_out0 = v$RM_3559_out0;
assign v$RM_11727_out0 = v$RM_3560_out0;
assign v$RM_11729_out0 = v$RM_3561_out0;
assign v$RM_11731_out0 = v$RM_3562_out0;
assign v$RM_11733_out0 = v$RM_3563_out0;
assign v$RM_12168_out0 = v$RM_3773_out0;
assign v$RM_12170_out0 = v$RM_3774_out0;
assign v$RM_12174_out0 = v$RM_3776_out0;
assign v$RM_12176_out0 = v$RM_3777_out0;
assign v$RM_12178_out0 = v$RM_3778_out0;
assign v$RM_12181_out0 = v$RM_3779_out0;
assign v$RM_12183_out0 = v$RM_3780_out0;
assign v$RM_12185_out0 = v$RM_3781_out0;
assign v$RM_12187_out0 = v$RM_3782_out0;
assign v$RM_12189_out0 = v$RM_3783_out0;
assign v$RM_12191_out0 = v$RM_3784_out0;
assign v$RM_12193_out0 = v$RM_3785_out0;
assign v$RM_12195_out0 = v$RM_3786_out0;
assign v$RM_12197_out0 = v$RM_3787_out0;
assign v$G2_12667_out0 = v$RD_6276_out0 && v$RM_11716_out0;
assign v$G2_13131_out0 = v$RD_6740_out0 && v$RM_12180_out0;
assign v$CARRY_5276_out0 = v$G2_12667_out0;
assign v$CARRY_5740_out0 = v$G2_13131_out0;
assign v$G1_8119_out0 = ((v$RD_6264_out0 && !v$RM_11704_out0) || (!v$RD_6264_out0) && v$RM_11704_out0);
assign v$G1_8121_out0 = ((v$RD_6266_out0 && !v$RM_11706_out0) || (!v$RD_6266_out0) && v$RM_11706_out0);
assign v$G1_8125_out0 = ((v$RD_6270_out0 && !v$RM_11710_out0) || (!v$RD_6270_out0) && v$RM_11710_out0);
assign v$G1_8127_out0 = ((v$RD_6272_out0 && !v$RM_11712_out0) || (!v$RD_6272_out0) && v$RM_11712_out0);
assign v$G1_8129_out0 = ((v$RD_6274_out0 && !v$RM_11714_out0) || (!v$RD_6274_out0) && v$RM_11714_out0);
assign v$G1_8132_out0 = ((v$RD_6277_out0 && !v$RM_11717_out0) || (!v$RD_6277_out0) && v$RM_11717_out0);
assign v$G1_8134_out0 = ((v$RD_6279_out0 && !v$RM_11719_out0) || (!v$RD_6279_out0) && v$RM_11719_out0);
assign v$G1_8136_out0 = ((v$RD_6281_out0 && !v$RM_11721_out0) || (!v$RD_6281_out0) && v$RM_11721_out0);
assign v$G1_8138_out0 = ((v$RD_6283_out0 && !v$RM_11723_out0) || (!v$RD_6283_out0) && v$RM_11723_out0);
assign v$G1_8140_out0 = ((v$RD_6285_out0 && !v$RM_11725_out0) || (!v$RD_6285_out0) && v$RM_11725_out0);
assign v$G1_8142_out0 = ((v$RD_6287_out0 && !v$RM_11727_out0) || (!v$RD_6287_out0) && v$RM_11727_out0);
assign v$G1_8144_out0 = ((v$RD_6289_out0 && !v$RM_11729_out0) || (!v$RD_6289_out0) && v$RM_11729_out0);
assign v$G1_8146_out0 = ((v$RD_6291_out0 && !v$RM_11731_out0) || (!v$RD_6291_out0) && v$RM_11731_out0);
assign v$G1_8148_out0 = ((v$RD_6293_out0 && !v$RM_11733_out0) || (!v$RD_6293_out0) && v$RM_11733_out0);
assign v$G1_8583_out0 = ((v$RD_6728_out0 && !v$RM_12168_out0) || (!v$RD_6728_out0) && v$RM_12168_out0);
assign v$G1_8585_out0 = ((v$RD_6730_out0 && !v$RM_12170_out0) || (!v$RD_6730_out0) && v$RM_12170_out0);
assign v$G1_8589_out0 = ((v$RD_6734_out0 && !v$RM_12174_out0) || (!v$RD_6734_out0) && v$RM_12174_out0);
assign v$G1_8591_out0 = ((v$RD_6736_out0 && !v$RM_12176_out0) || (!v$RD_6736_out0) && v$RM_12176_out0);
assign v$G1_8593_out0 = ((v$RD_6738_out0 && !v$RM_12178_out0) || (!v$RD_6738_out0) && v$RM_12178_out0);
assign v$G1_8596_out0 = ((v$RD_6741_out0 && !v$RM_12181_out0) || (!v$RD_6741_out0) && v$RM_12181_out0);
assign v$G1_8598_out0 = ((v$RD_6743_out0 && !v$RM_12183_out0) || (!v$RD_6743_out0) && v$RM_12183_out0);
assign v$G1_8600_out0 = ((v$RD_6745_out0 && !v$RM_12185_out0) || (!v$RD_6745_out0) && v$RM_12185_out0);
assign v$G1_8602_out0 = ((v$RD_6747_out0 && !v$RM_12187_out0) || (!v$RD_6747_out0) && v$RM_12187_out0);
assign v$G1_8604_out0 = ((v$RD_6749_out0 && !v$RM_12189_out0) || (!v$RD_6749_out0) && v$RM_12189_out0);
assign v$G1_8606_out0 = ((v$RD_6751_out0 && !v$RM_12191_out0) || (!v$RD_6751_out0) && v$RM_12191_out0);
assign v$G1_8608_out0 = ((v$RD_6753_out0 && !v$RM_12193_out0) || (!v$RD_6753_out0) && v$RM_12193_out0);
assign v$G1_8610_out0 = ((v$RD_6755_out0 && !v$RM_12195_out0) || (!v$RD_6755_out0) && v$RM_12195_out0);
assign v$G1_8612_out0 = ((v$RD_6757_out0 && !v$RM_12197_out0) || (!v$RD_6757_out0) && v$RM_12197_out0);
assign v$S_9277_out0 = v$G1_8131_out0;
assign v$S_9741_out0 = v$G1_8595_out0;
assign v$G2_12655_out0 = v$RD_6264_out0 && v$RM_11704_out0;
assign v$G2_12657_out0 = v$RD_6266_out0 && v$RM_11706_out0;
assign v$G2_12661_out0 = v$RD_6270_out0 && v$RM_11710_out0;
assign v$G2_12663_out0 = v$RD_6272_out0 && v$RM_11712_out0;
assign v$G2_12665_out0 = v$RD_6274_out0 && v$RM_11714_out0;
assign v$G2_12668_out0 = v$RD_6277_out0 && v$RM_11717_out0;
assign v$G2_12670_out0 = v$RD_6279_out0 && v$RM_11719_out0;
assign v$G2_12672_out0 = v$RD_6281_out0 && v$RM_11721_out0;
assign v$G2_12674_out0 = v$RD_6283_out0 && v$RM_11723_out0;
assign v$G2_12676_out0 = v$RD_6285_out0 && v$RM_11725_out0;
assign v$G2_12678_out0 = v$RD_6287_out0 && v$RM_11727_out0;
assign v$G2_12680_out0 = v$RD_6289_out0 && v$RM_11729_out0;
assign v$G2_12682_out0 = v$RD_6291_out0 && v$RM_11731_out0;
assign v$G2_12684_out0 = v$RD_6293_out0 && v$RM_11733_out0;
assign v$G2_13119_out0 = v$RD_6728_out0 && v$RM_12168_out0;
assign v$G2_13121_out0 = v$RD_6730_out0 && v$RM_12170_out0;
assign v$G2_13125_out0 = v$RD_6734_out0 && v$RM_12174_out0;
assign v$G2_13127_out0 = v$RD_6736_out0 && v$RM_12176_out0;
assign v$G2_13129_out0 = v$RD_6738_out0 && v$RM_12178_out0;
assign v$G2_13132_out0 = v$RD_6741_out0 && v$RM_12181_out0;
assign v$G2_13134_out0 = v$RD_6743_out0 && v$RM_12183_out0;
assign v$G2_13136_out0 = v$RD_6745_out0 && v$RM_12185_out0;
assign v$G2_13138_out0 = v$RD_6747_out0 && v$RM_12187_out0;
assign v$G2_13140_out0 = v$RD_6749_out0 && v$RM_12189_out0;
assign v$G2_13142_out0 = v$RD_6751_out0 && v$RM_12191_out0;
assign v$G2_13144_out0 = v$RD_6753_out0 && v$RM_12193_out0;
assign v$G2_13146_out0 = v$RD_6755_out0 && v$RM_12195_out0;
assign v$G2_13148_out0 = v$RD_6757_out0 && v$RM_12197_out0;
assign v$S_4678_out0 = v$S_9277_out0;
assign v$S_4693_out0 = v$S_9741_out0;
assign v$CARRY_5264_out0 = v$G2_12655_out0;
assign v$CARRY_5266_out0 = v$G2_12657_out0;
assign v$CARRY_5270_out0 = v$G2_12661_out0;
assign v$CARRY_5272_out0 = v$G2_12663_out0;
assign v$CARRY_5274_out0 = v$G2_12665_out0;
assign v$CARRY_5277_out0 = v$G2_12668_out0;
assign v$CARRY_5279_out0 = v$G2_12670_out0;
assign v$CARRY_5281_out0 = v$G2_12672_out0;
assign v$CARRY_5283_out0 = v$G2_12674_out0;
assign v$CARRY_5285_out0 = v$G2_12676_out0;
assign v$CARRY_5287_out0 = v$G2_12678_out0;
assign v$CARRY_5289_out0 = v$G2_12680_out0;
assign v$CARRY_5291_out0 = v$G2_12682_out0;
assign v$CARRY_5293_out0 = v$G2_12684_out0;
assign v$CARRY_5728_out0 = v$G2_13119_out0;
assign v$CARRY_5730_out0 = v$G2_13121_out0;
assign v$CARRY_5734_out0 = v$G2_13125_out0;
assign v$CARRY_5736_out0 = v$G2_13127_out0;
assign v$CARRY_5738_out0 = v$G2_13129_out0;
assign v$CARRY_5741_out0 = v$G2_13132_out0;
assign v$CARRY_5743_out0 = v$G2_13134_out0;
assign v$CARRY_5745_out0 = v$G2_13136_out0;
assign v$CARRY_5747_out0 = v$G2_13138_out0;
assign v$CARRY_5749_out0 = v$G2_13140_out0;
assign v$CARRY_5751_out0 = v$G2_13142_out0;
assign v$CARRY_5753_out0 = v$G2_13144_out0;
assign v$CARRY_5755_out0 = v$G2_13146_out0;
assign v$CARRY_5757_out0 = v$G2_13148_out0;
assign v$S_9265_out0 = v$G1_8119_out0;
assign v$S_9267_out0 = v$G1_8121_out0;
assign v$S_9271_out0 = v$G1_8125_out0;
assign v$S_9273_out0 = v$G1_8127_out0;
assign v$S_9275_out0 = v$G1_8129_out0;
assign v$S_9278_out0 = v$G1_8132_out0;
assign v$S_9280_out0 = v$G1_8134_out0;
assign v$S_9282_out0 = v$G1_8136_out0;
assign v$S_9284_out0 = v$G1_8138_out0;
assign v$S_9286_out0 = v$G1_8140_out0;
assign v$S_9288_out0 = v$G1_8142_out0;
assign v$S_9290_out0 = v$G1_8144_out0;
assign v$S_9292_out0 = v$G1_8146_out0;
assign v$S_9294_out0 = v$G1_8148_out0;
assign v$S_9729_out0 = v$G1_8583_out0;
assign v$S_9731_out0 = v$G1_8585_out0;
assign v$S_9735_out0 = v$G1_8589_out0;
assign v$S_9737_out0 = v$G1_8591_out0;
assign v$S_9739_out0 = v$G1_8593_out0;
assign v$S_9742_out0 = v$G1_8596_out0;
assign v$S_9744_out0 = v$G1_8598_out0;
assign v$S_9746_out0 = v$G1_8600_out0;
assign v$S_9748_out0 = v$G1_8602_out0;
assign v$S_9750_out0 = v$G1_8604_out0;
assign v$S_9752_out0 = v$G1_8606_out0;
assign v$S_9754_out0 = v$G1_8608_out0;
assign v$S_9756_out0 = v$G1_8610_out0;
assign v$S_9758_out0 = v$G1_8612_out0;
assign v$CIN_10010_out0 = v$CARRY_5276_out0;
assign v$CIN_10234_out0 = v$CARRY_5740_out0;
assign v$_681_out0 = { v$_56_out0,v$S_4678_out0 };
assign v$_682_out0 = { v$_57_out0,v$S_4693_out0 };
assign v$RD_6282_out0 = v$CIN_10010_out0;
assign v$RD_6746_out0 = v$CIN_10234_out0;
assign v$RM_11705_out0 = v$S_9265_out0;
assign v$RM_11707_out0 = v$S_9267_out0;
assign v$RM_11711_out0 = v$S_9271_out0;
assign v$RM_11713_out0 = v$S_9273_out0;
assign v$RM_11715_out0 = v$S_9275_out0;
assign v$RM_11718_out0 = v$S_9278_out0;
assign v$RM_11720_out0 = v$S_9280_out0;
assign v$RM_11722_out0 = v$S_9282_out0;
assign v$RM_11724_out0 = v$S_9284_out0;
assign v$RM_11726_out0 = v$S_9286_out0;
assign v$RM_11728_out0 = v$S_9288_out0;
assign v$RM_11730_out0 = v$S_9290_out0;
assign v$RM_11732_out0 = v$S_9292_out0;
assign v$RM_11734_out0 = v$S_9294_out0;
assign v$RM_12169_out0 = v$S_9729_out0;
assign v$RM_12171_out0 = v$S_9731_out0;
assign v$RM_12175_out0 = v$S_9735_out0;
assign v$RM_12177_out0 = v$S_9737_out0;
assign v$RM_12179_out0 = v$S_9739_out0;
assign v$RM_12182_out0 = v$S_9742_out0;
assign v$RM_12184_out0 = v$S_9744_out0;
assign v$RM_12186_out0 = v$S_9746_out0;
assign v$RM_12188_out0 = v$S_9748_out0;
assign v$RM_12190_out0 = v$S_9750_out0;
assign v$RM_12192_out0 = v$S_9752_out0;
assign v$RM_12194_out0 = v$S_9754_out0;
assign v$RM_12196_out0 = v$S_9756_out0;
assign v$RM_12198_out0 = v$S_9758_out0;
assign v$G1_8137_out0 = ((v$RD_6282_out0 && !v$RM_11722_out0) || (!v$RD_6282_out0) && v$RM_11722_out0);
assign v$G1_8601_out0 = ((v$RD_6746_out0 && !v$RM_12186_out0) || (!v$RD_6746_out0) && v$RM_12186_out0);
assign v$G2_12673_out0 = v$RD_6282_out0 && v$RM_11722_out0;
assign v$G2_13137_out0 = v$RD_6746_out0 && v$RM_12186_out0;
assign v$CARRY_5282_out0 = v$G2_12673_out0;
assign v$CARRY_5746_out0 = v$G2_13137_out0;
assign v$S_9283_out0 = v$G1_8137_out0;
assign v$S_9747_out0 = v$G1_8601_out0;
assign v$S_1421_out0 = v$S_9283_out0;
assign v$S_1645_out0 = v$S_9747_out0;
assign v$G1_4197_out0 = v$CARRY_5282_out0 || v$CARRY_5281_out0;
assign v$G1_4421_out0 = v$CARRY_5746_out0 || v$CARRY_5745_out0;
assign v$COUT_889_out0 = v$G1_4197_out0;
assign v$COUT_1113_out0 = v$G1_4421_out0;
assign v$CIN_10016_out0 = v$COUT_889_out0;
assign v$CIN_10240_out0 = v$COUT_1113_out0;
assign v$RD_6294_out0 = v$CIN_10016_out0;
assign v$RD_6758_out0 = v$CIN_10240_out0;
assign v$G1_8149_out0 = ((v$RD_6294_out0 && !v$RM_11734_out0) || (!v$RD_6294_out0) && v$RM_11734_out0);
assign v$G1_8613_out0 = ((v$RD_6758_out0 && !v$RM_12198_out0) || (!v$RD_6758_out0) && v$RM_12198_out0);
assign v$G2_12685_out0 = v$RD_6294_out0 && v$RM_11734_out0;
assign v$G2_13149_out0 = v$RD_6758_out0 && v$RM_12198_out0;
assign v$CARRY_5294_out0 = v$G2_12685_out0;
assign v$CARRY_5758_out0 = v$G2_13149_out0;
assign v$S_9295_out0 = v$G1_8149_out0;
assign v$S_9759_out0 = v$G1_8613_out0;
assign v$S_1427_out0 = v$S_9295_out0;
assign v$S_1651_out0 = v$S_9759_out0;
assign v$G1_4203_out0 = v$CARRY_5294_out0 || v$CARRY_5293_out0;
assign v$G1_4427_out0 = v$CARRY_5758_out0 || v$CARRY_5757_out0;
assign v$COUT_895_out0 = v$G1_4203_out0;
assign v$COUT_1119_out0 = v$G1_4427_out0;
assign v$_4795_out0 = { v$S_1421_out0,v$S_1427_out0 };
assign v$_4810_out0 = { v$S_1645_out0,v$S_1651_out0 };
assign v$CIN_10011_out0 = v$COUT_895_out0;
assign v$CIN_10235_out0 = v$COUT_1119_out0;
assign v$RD_6284_out0 = v$CIN_10011_out0;
assign v$RD_6748_out0 = v$CIN_10235_out0;
assign v$G1_8139_out0 = ((v$RD_6284_out0 && !v$RM_11724_out0) || (!v$RD_6284_out0) && v$RM_11724_out0);
assign v$G1_8603_out0 = ((v$RD_6748_out0 && !v$RM_12188_out0) || (!v$RD_6748_out0) && v$RM_12188_out0);
assign v$G2_12675_out0 = v$RD_6284_out0 && v$RM_11724_out0;
assign v$G2_13139_out0 = v$RD_6748_out0 && v$RM_12188_out0;
assign v$CARRY_5284_out0 = v$G2_12675_out0;
assign v$CARRY_5748_out0 = v$G2_13139_out0;
assign v$S_9285_out0 = v$G1_8139_out0;
assign v$S_9749_out0 = v$G1_8603_out0;
assign v$S_1422_out0 = v$S_9285_out0;
assign v$S_1646_out0 = v$S_9749_out0;
assign v$G1_4198_out0 = v$CARRY_5284_out0 || v$CARRY_5283_out0;
assign v$G1_4422_out0 = v$CARRY_5748_out0 || v$CARRY_5747_out0;
assign v$COUT_890_out0 = v$G1_4198_out0;
assign v$COUT_1114_out0 = v$G1_4422_out0;
assign v$_2565_out0 = { v$_4795_out0,v$S_1422_out0 };
assign v$_2580_out0 = { v$_4810_out0,v$S_1646_out0 };
assign v$CIN_10006_out0 = v$COUT_890_out0;
assign v$CIN_10230_out0 = v$COUT_1114_out0;
assign v$RD_6273_out0 = v$CIN_10006_out0;
assign v$RD_6737_out0 = v$CIN_10230_out0;
assign v$G1_8128_out0 = ((v$RD_6273_out0 && !v$RM_11713_out0) || (!v$RD_6273_out0) && v$RM_11713_out0);
assign v$G1_8592_out0 = ((v$RD_6737_out0 && !v$RM_12177_out0) || (!v$RD_6737_out0) && v$RM_12177_out0);
assign v$G2_12664_out0 = v$RD_6273_out0 && v$RM_11713_out0;
assign v$G2_13128_out0 = v$RD_6737_out0 && v$RM_12177_out0;
assign v$CARRY_5273_out0 = v$G2_12664_out0;
assign v$CARRY_5737_out0 = v$G2_13128_out0;
assign v$S_9274_out0 = v$G1_8128_out0;
assign v$S_9738_out0 = v$G1_8592_out0;
assign v$S_1417_out0 = v$S_9274_out0;
assign v$S_1641_out0 = v$S_9738_out0;
assign v$G1_4193_out0 = v$CARRY_5273_out0 || v$CARRY_5272_out0;
assign v$G1_4417_out0 = v$CARRY_5737_out0 || v$CARRY_5736_out0;
assign v$COUT_885_out0 = v$G1_4193_out0;
assign v$COUT_1109_out0 = v$G1_4417_out0;
assign v$_7045_out0 = { v$_2565_out0,v$S_1417_out0 };
assign v$_7060_out0 = { v$_2580_out0,v$S_1641_out0 };
assign v$CIN_10005_out0 = v$COUT_885_out0;
assign v$CIN_10229_out0 = v$COUT_1109_out0;
assign v$RD_6271_out0 = v$CIN_10005_out0;
assign v$RD_6735_out0 = v$CIN_10229_out0;
assign v$G1_8126_out0 = ((v$RD_6271_out0 && !v$RM_11711_out0) || (!v$RD_6271_out0) && v$RM_11711_out0);
assign v$G1_8590_out0 = ((v$RD_6735_out0 && !v$RM_12175_out0) || (!v$RD_6735_out0) && v$RM_12175_out0);
assign v$G2_12662_out0 = v$RD_6271_out0 && v$RM_11711_out0;
assign v$G2_13126_out0 = v$RD_6735_out0 && v$RM_12175_out0;
assign v$CARRY_5271_out0 = v$G2_12662_out0;
assign v$CARRY_5735_out0 = v$G2_13126_out0;
assign v$S_9272_out0 = v$G1_8126_out0;
assign v$S_9736_out0 = v$G1_8590_out0;
assign v$S_1416_out0 = v$S_9272_out0;
assign v$S_1640_out0 = v$S_9736_out0;
assign v$G1_4192_out0 = v$CARRY_5271_out0 || v$CARRY_5270_out0;
assign v$G1_4416_out0 = v$CARRY_5735_out0 || v$CARRY_5734_out0;
assign v$COUT_884_out0 = v$G1_4192_out0;
assign v$COUT_1108_out0 = v$G1_4416_out0;
assign v$_13531_out0 = { v$_7045_out0,v$S_1416_out0 };
assign v$_13546_out0 = { v$_7060_out0,v$S_1640_out0 };
assign v$CIN_10012_out0 = v$COUT_884_out0;
assign v$CIN_10236_out0 = v$COUT_1108_out0;
assign v$RD_6286_out0 = v$CIN_10012_out0;
assign v$RD_6750_out0 = v$CIN_10236_out0;
assign v$G1_8141_out0 = ((v$RD_6286_out0 && !v$RM_11726_out0) || (!v$RD_6286_out0) && v$RM_11726_out0);
assign v$G1_8605_out0 = ((v$RD_6750_out0 && !v$RM_12190_out0) || (!v$RD_6750_out0) && v$RM_12190_out0);
assign v$G2_12677_out0 = v$RD_6286_out0 && v$RM_11726_out0;
assign v$G2_13141_out0 = v$RD_6750_out0 && v$RM_12190_out0;
assign v$CARRY_5286_out0 = v$G2_12677_out0;
assign v$CARRY_5750_out0 = v$G2_13141_out0;
assign v$S_9287_out0 = v$G1_8141_out0;
assign v$S_9751_out0 = v$G1_8605_out0;
assign v$S_1423_out0 = v$S_9287_out0;
assign v$S_1647_out0 = v$S_9751_out0;
assign v$G1_4199_out0 = v$CARRY_5286_out0 || v$CARRY_5285_out0;
assign v$G1_4423_out0 = v$CARRY_5750_out0 || v$CARRY_5749_out0;
assign v$COUT_891_out0 = v$G1_4199_out0;
assign v$COUT_1115_out0 = v$G1_4423_out0;
assign v$_3324_out0 = { v$_13531_out0,v$S_1423_out0 };
assign v$_3339_out0 = { v$_13546_out0,v$S_1647_out0 };
assign v$CIN_10013_out0 = v$COUT_891_out0;
assign v$CIN_10237_out0 = v$COUT_1115_out0;
assign v$RD_6288_out0 = v$CIN_10013_out0;
assign v$RD_6752_out0 = v$CIN_10237_out0;
assign v$G1_8143_out0 = ((v$RD_6288_out0 && !v$RM_11728_out0) || (!v$RD_6288_out0) && v$RM_11728_out0);
assign v$G1_8607_out0 = ((v$RD_6752_out0 && !v$RM_12192_out0) || (!v$RD_6752_out0) && v$RM_12192_out0);
assign v$G2_12679_out0 = v$RD_6288_out0 && v$RM_11728_out0;
assign v$G2_13143_out0 = v$RD_6752_out0 && v$RM_12192_out0;
assign v$CARRY_5288_out0 = v$G2_12679_out0;
assign v$CARRY_5752_out0 = v$G2_13143_out0;
assign v$S_9289_out0 = v$G1_8143_out0;
assign v$S_9753_out0 = v$G1_8607_out0;
assign v$S_1424_out0 = v$S_9289_out0;
assign v$S_1648_out0 = v$S_9753_out0;
assign v$G1_4200_out0 = v$CARRY_5288_out0 || v$CARRY_5287_out0;
assign v$G1_4424_out0 = v$CARRY_5752_out0 || v$CARRY_5751_out0;
assign v$COUT_892_out0 = v$G1_4200_out0;
assign v$COUT_1116_out0 = v$G1_4424_out0;
assign v$_7160_out0 = { v$_3324_out0,v$S_1424_out0 };
assign v$_7175_out0 = { v$_3339_out0,v$S_1648_out0 };
assign v$CIN_10015_out0 = v$COUT_892_out0;
assign v$CIN_10239_out0 = v$COUT_1116_out0;
assign v$RD_6292_out0 = v$CIN_10015_out0;
assign v$RD_6756_out0 = v$CIN_10239_out0;
assign v$G1_8147_out0 = ((v$RD_6292_out0 && !v$RM_11732_out0) || (!v$RD_6292_out0) && v$RM_11732_out0);
assign v$G1_8611_out0 = ((v$RD_6756_out0 && !v$RM_12196_out0) || (!v$RD_6756_out0) && v$RM_12196_out0);
assign v$G2_12683_out0 = v$RD_6292_out0 && v$RM_11732_out0;
assign v$G2_13147_out0 = v$RD_6756_out0 && v$RM_12196_out0;
assign v$CARRY_5292_out0 = v$G2_12683_out0;
assign v$CARRY_5756_out0 = v$G2_13147_out0;
assign v$S_9293_out0 = v$G1_8147_out0;
assign v$S_9757_out0 = v$G1_8611_out0;
assign v$S_1426_out0 = v$S_9293_out0;
assign v$S_1650_out0 = v$S_9757_out0;
assign v$G1_4202_out0 = v$CARRY_5292_out0 || v$CARRY_5291_out0;
assign v$G1_4426_out0 = v$CARRY_5756_out0 || v$CARRY_5755_out0;
assign v$COUT_894_out0 = v$G1_4202_out0;
assign v$COUT_1118_out0 = v$G1_4426_out0;
assign v$_4762_out0 = { v$_7160_out0,v$S_1426_out0 };
assign v$_4777_out0 = { v$_7175_out0,v$S_1650_out0 };
assign v$CIN_10008_out0 = v$COUT_894_out0;
assign v$CIN_10232_out0 = v$COUT_1118_out0;
assign v$RD_6278_out0 = v$CIN_10008_out0;
assign v$RD_6742_out0 = v$CIN_10232_out0;
assign v$G1_8133_out0 = ((v$RD_6278_out0 && !v$RM_11718_out0) || (!v$RD_6278_out0) && v$RM_11718_out0);
assign v$G1_8597_out0 = ((v$RD_6742_out0 && !v$RM_12182_out0) || (!v$RD_6742_out0) && v$RM_12182_out0);
assign v$G2_12669_out0 = v$RD_6278_out0 && v$RM_11718_out0;
assign v$G2_13133_out0 = v$RD_6742_out0 && v$RM_12182_out0;
assign v$CARRY_5278_out0 = v$G2_12669_out0;
assign v$CARRY_5742_out0 = v$G2_13133_out0;
assign v$S_9279_out0 = v$G1_8133_out0;
assign v$S_9743_out0 = v$G1_8597_out0;
assign v$S_1419_out0 = v$S_9279_out0;
assign v$S_1643_out0 = v$S_9743_out0;
assign v$G1_4195_out0 = v$CARRY_5278_out0 || v$CARRY_5277_out0;
assign v$G1_4419_out0 = v$CARRY_5742_out0 || v$CARRY_5741_out0;
assign v$COUT_887_out0 = v$G1_4195_out0;
assign v$COUT_1111_out0 = v$G1_4419_out0;
assign v$_6939_out0 = { v$_4762_out0,v$S_1419_out0 };
assign v$_6954_out0 = { v$_4777_out0,v$S_1643_out0 };
assign v$CIN_10009_out0 = v$COUT_887_out0;
assign v$CIN_10233_out0 = v$COUT_1111_out0;
assign v$RD_6280_out0 = v$CIN_10009_out0;
assign v$RD_6744_out0 = v$CIN_10233_out0;
assign v$G1_8135_out0 = ((v$RD_6280_out0 && !v$RM_11720_out0) || (!v$RD_6280_out0) && v$RM_11720_out0);
assign v$G1_8599_out0 = ((v$RD_6744_out0 && !v$RM_12184_out0) || (!v$RD_6744_out0) && v$RM_12184_out0);
assign v$G2_12671_out0 = v$RD_6280_out0 && v$RM_11720_out0;
assign v$G2_13135_out0 = v$RD_6744_out0 && v$RM_12184_out0;
assign v$CARRY_5280_out0 = v$G2_12671_out0;
assign v$CARRY_5744_out0 = v$G2_13135_out0;
assign v$S_9281_out0 = v$G1_8135_out0;
assign v$S_9745_out0 = v$G1_8599_out0;
assign v$S_1420_out0 = v$S_9281_out0;
assign v$S_1644_out0 = v$S_9745_out0;
assign v$G1_4196_out0 = v$CARRY_5280_out0 || v$CARRY_5279_out0;
assign v$G1_4420_out0 = v$CARRY_5744_out0 || v$CARRY_5743_out0;
assign v$COUT_888_out0 = v$G1_4196_out0;
assign v$COUT_1112_out0 = v$G1_4420_out0;
assign v$_5815_out0 = { v$_6939_out0,v$S_1420_out0 };
assign v$_5830_out0 = { v$_6954_out0,v$S_1644_out0 };
assign v$CIN_10014_out0 = v$COUT_888_out0;
assign v$CIN_10238_out0 = v$COUT_1112_out0;
assign v$RD_6290_out0 = v$CIN_10014_out0;
assign v$RD_6754_out0 = v$CIN_10238_out0;
assign v$G1_8145_out0 = ((v$RD_6290_out0 && !v$RM_11730_out0) || (!v$RD_6290_out0) && v$RM_11730_out0);
assign v$G1_8609_out0 = ((v$RD_6754_out0 && !v$RM_12194_out0) || (!v$RD_6754_out0) && v$RM_12194_out0);
assign v$G2_12681_out0 = v$RD_6290_out0 && v$RM_11730_out0;
assign v$G2_13145_out0 = v$RD_6754_out0 && v$RM_12194_out0;
assign v$CARRY_5290_out0 = v$G2_12681_out0;
assign v$CARRY_5754_out0 = v$G2_13145_out0;
assign v$S_9291_out0 = v$G1_8145_out0;
assign v$S_9755_out0 = v$G1_8609_out0;
assign v$S_1425_out0 = v$S_9291_out0;
assign v$S_1649_out0 = v$S_9755_out0;
assign v$G1_4201_out0 = v$CARRY_5290_out0 || v$CARRY_5289_out0;
assign v$G1_4425_out0 = v$CARRY_5754_out0 || v$CARRY_5753_out0;
assign v$COUT_893_out0 = v$G1_4201_out0;
assign v$COUT_1117_out0 = v$G1_4425_out0;
assign v$_2039_out0 = { v$_5815_out0,v$S_1425_out0 };
assign v$_2054_out0 = { v$_5830_out0,v$S_1649_out0 };
assign v$CIN_10002_out0 = v$COUT_893_out0;
assign v$CIN_10226_out0 = v$COUT_1117_out0;
assign v$RD_6265_out0 = v$CIN_10002_out0;
assign v$RD_6729_out0 = v$CIN_10226_out0;
assign v$G1_8120_out0 = ((v$RD_6265_out0 && !v$RM_11705_out0) || (!v$RD_6265_out0) && v$RM_11705_out0);
assign v$G1_8584_out0 = ((v$RD_6729_out0 && !v$RM_12169_out0) || (!v$RD_6729_out0) && v$RM_12169_out0);
assign v$G2_12656_out0 = v$RD_6265_out0 && v$RM_11705_out0;
assign v$G2_13120_out0 = v$RD_6729_out0 && v$RM_12169_out0;
assign v$CARRY_5265_out0 = v$G2_12656_out0;
assign v$CARRY_5729_out0 = v$G2_13120_out0;
assign v$S_9266_out0 = v$G1_8120_out0;
assign v$S_9730_out0 = v$G1_8584_out0;
assign v$S_1413_out0 = v$S_9266_out0;
assign v$S_1637_out0 = v$S_9730_out0;
assign v$G1_4189_out0 = v$CARRY_5265_out0 || v$CARRY_5264_out0;
assign v$G1_4413_out0 = v$CARRY_5729_out0 || v$CARRY_5728_out0;
assign v$COUT_881_out0 = v$G1_4189_out0;
assign v$COUT_1105_out0 = v$G1_4413_out0;
assign v$_2806_out0 = { v$_2039_out0,v$S_1413_out0 };
assign v$_2821_out0 = { v$_2054_out0,v$S_1637_out0 };
assign v$CIN_10007_out0 = v$COUT_881_out0;
assign v$CIN_10231_out0 = v$COUT_1105_out0;
assign v$RD_6275_out0 = v$CIN_10007_out0;
assign v$RD_6739_out0 = v$CIN_10231_out0;
assign v$G1_8130_out0 = ((v$RD_6275_out0 && !v$RM_11715_out0) || (!v$RD_6275_out0) && v$RM_11715_out0);
assign v$G1_8594_out0 = ((v$RD_6739_out0 && !v$RM_12179_out0) || (!v$RD_6739_out0) && v$RM_12179_out0);
assign v$G2_12666_out0 = v$RD_6275_out0 && v$RM_11715_out0;
assign v$G2_13130_out0 = v$RD_6739_out0 && v$RM_12179_out0;
assign v$CARRY_5275_out0 = v$G2_12666_out0;
assign v$CARRY_5739_out0 = v$G2_13130_out0;
assign v$S_9276_out0 = v$G1_8130_out0;
assign v$S_9740_out0 = v$G1_8594_out0;
assign v$S_1418_out0 = v$S_9276_out0;
assign v$S_1642_out0 = v$S_9740_out0;
assign v$G1_4194_out0 = v$CARRY_5275_out0 || v$CARRY_5274_out0;
assign v$G1_4418_out0 = v$CARRY_5739_out0 || v$CARRY_5738_out0;
assign v$COUT_886_out0 = v$G1_4194_out0;
assign v$COUT_1110_out0 = v$G1_4418_out0;
assign v$_1838_out0 = { v$_2806_out0,v$S_1418_out0 };
assign v$_1853_out0 = { v$_2821_out0,v$S_1642_out0 };
assign v$CIN_10003_out0 = v$COUT_886_out0;
assign v$CIN_10227_out0 = v$COUT_1110_out0;
assign v$RD_6267_out0 = v$CIN_10003_out0;
assign v$RD_6731_out0 = v$CIN_10227_out0;
assign v$G1_8122_out0 = ((v$RD_6267_out0 && !v$RM_11707_out0) || (!v$RD_6267_out0) && v$RM_11707_out0);
assign v$G1_8586_out0 = ((v$RD_6731_out0 && !v$RM_12171_out0) || (!v$RD_6731_out0) && v$RM_12171_out0);
assign v$G2_12658_out0 = v$RD_6267_out0 && v$RM_11707_out0;
assign v$G2_13122_out0 = v$RD_6731_out0 && v$RM_12171_out0;
assign v$CARRY_5267_out0 = v$G2_12658_out0;
assign v$CARRY_5731_out0 = v$G2_13122_out0;
assign v$S_9268_out0 = v$G1_8122_out0;
assign v$S_9732_out0 = v$G1_8586_out0;
assign v$S_1414_out0 = v$S_9268_out0;
assign v$S_1638_out0 = v$S_9732_out0;
assign v$G1_4190_out0 = v$CARRY_5267_out0 || v$CARRY_5266_out0;
assign v$G1_4414_out0 = v$CARRY_5731_out0 || v$CARRY_5730_out0;
assign v$COUT_882_out0 = v$G1_4190_out0;
assign v$COUT_1106_out0 = v$G1_4414_out0;
assign v$_4562_out0 = { v$_1838_out0,v$S_1414_out0 };
assign v$_4577_out0 = { v$_1853_out0,v$S_1638_out0 };
assign v$RM_3551_out0 = v$COUT_882_out0;
assign v$RM_3775_out0 = v$COUT_1106_out0;
assign v$RM_11708_out0 = v$RM_3551_out0;
assign v$RM_12172_out0 = v$RM_3775_out0;
assign v$G1_8123_out0 = ((v$RD_6268_out0 && !v$RM_11708_out0) || (!v$RD_6268_out0) && v$RM_11708_out0);
assign v$G1_8587_out0 = ((v$RD_6732_out0 && !v$RM_12172_out0) || (!v$RD_6732_out0) && v$RM_12172_out0);
assign v$G2_12659_out0 = v$RD_6268_out0 && v$RM_11708_out0;
assign v$G2_13123_out0 = v$RD_6732_out0 && v$RM_12172_out0;
assign v$CARRY_5268_out0 = v$G2_12659_out0;
assign v$CARRY_5732_out0 = v$G2_13123_out0;
assign v$S_9269_out0 = v$G1_8123_out0;
assign v$S_9733_out0 = v$G1_8587_out0;
assign v$RM_11709_out0 = v$S_9269_out0;
assign v$RM_12173_out0 = v$S_9733_out0;
assign v$G1_8124_out0 = ((v$RD_6269_out0 && !v$RM_11709_out0) || (!v$RD_6269_out0) && v$RM_11709_out0);
assign v$G1_8588_out0 = ((v$RD_6733_out0 && !v$RM_12173_out0) || (!v$RD_6733_out0) && v$RM_12173_out0);
assign v$G2_12660_out0 = v$RD_6269_out0 && v$RM_11709_out0;
assign v$G2_13124_out0 = v$RD_6733_out0 && v$RM_12173_out0;
assign v$CARRY_5269_out0 = v$G2_12660_out0;
assign v$CARRY_5733_out0 = v$G2_13124_out0;
assign v$S_9270_out0 = v$G1_8124_out0;
assign v$S_9734_out0 = v$G1_8588_out0;
assign v$S_1415_out0 = v$S_9270_out0;
assign v$S_1639_out0 = v$S_9734_out0;
assign v$G1_4191_out0 = v$CARRY_5269_out0 || v$CARRY_5268_out0;
assign v$G1_4415_out0 = v$CARRY_5733_out0 || v$CARRY_5732_out0;
assign v$COUT_883_out0 = v$G1_4191_out0;
assign v$COUT_1107_out0 = v$G1_4415_out0;
assign v$_10664_out0 = { v$_4562_out0,v$S_1415_out0 };
assign v$_10679_out0 = { v$_4577_out0,v$S_1639_out0 };
assign v$_10959_out0 = { v$_10664_out0,v$COUT_883_out0 };
assign v$_10974_out0 = { v$_10679_out0,v$COUT_1107_out0 };
assign v$COUT_10929_out0 = v$_10959_out0;
assign v$COUT_10944_out0 = v$_10974_out0;
assign v$CIN_2366_out0 = v$COUT_10929_out0;
assign v$CIN_2381_out0 = v$COUT_10944_out0;
assign v$_479_out0 = v$CIN_2366_out0[8:8];
assign v$_494_out0 = v$CIN_2381_out0[8:8];
assign v$_1784_out0 = v$CIN_2366_out0[6:6];
assign v$_1799_out0 = v$CIN_2381_out0[6:6];
assign v$_2166_out0 = v$CIN_2366_out0[3:3];
assign v$_2181_out0 = v$CIN_2381_out0[3:3];
assign v$_2205_out0 = v$CIN_2366_out0[15:15];
assign v$_2219_out0 = v$CIN_2381_out0[15:15];
assign v$_2513_out0 = v$CIN_2366_out0[0:0];
assign v$_2528_out0 = v$CIN_2381_out0[0:0];
assign v$_3062_out0 = v$CIN_2366_out0[9:9];
assign v$_3077_out0 = v$CIN_2381_out0[9:9];
assign v$_3096_out0 = v$CIN_2366_out0[2:2];
assign v$_3111_out0 = v$CIN_2381_out0[2:2];
assign v$_3150_out0 = v$CIN_2366_out0[7:7];
assign v$_3165_out0 = v$CIN_2381_out0[7:7];
assign v$_3834_out0 = v$CIN_2366_out0[1:1];
assign v$_3849_out0 = v$CIN_2381_out0[1:1];
assign v$_3872_out0 = v$CIN_2366_out0[10:10];
assign v$_3887_out0 = v$CIN_2381_out0[10:10];
assign v$_6811_out0 = v$CIN_2366_out0[11:11];
assign v$_6826_out0 = v$CIN_2381_out0[11:11];
assign v$_7655_out0 = v$CIN_2366_out0[12:12];
assign v$_7670_out0 = v$CIN_2381_out0[12:12];
assign v$_8710_out0 = v$CIN_2366_out0[13:13];
assign v$_8725_out0 = v$CIN_2381_out0[13:13];
assign v$_8780_out0 = v$CIN_2366_out0[14:14];
assign v$_8795_out0 = v$CIN_2381_out0[14:14];
assign v$_10730_out0 = v$CIN_2366_out0[5:5];
assign v$_10745_out0 = v$CIN_2381_out0[5:5];
assign v$_13459_out0 = v$CIN_2366_out0[4:4];
assign v$_13474_out0 = v$CIN_2381_out0[4:4];
assign v$RM_3519_out0 = v$_7655_out0;
assign v$RM_3520_out0 = v$_8780_out0;
assign v$RM_3522_out0 = v$_10730_out0;
assign v$RM_3523_out0 = v$_13459_out0;
assign v$RM_3524_out0 = v$_8710_out0;
assign v$RM_3525_out0 = v$_3062_out0;
assign v$RM_3526_out0 = v$_3872_out0;
assign v$RM_3527_out0 = v$_3834_out0;
assign v$RM_3528_out0 = v$_2166_out0;
assign v$RM_3529_out0 = v$_1784_out0;
assign v$RM_3530_out0 = v$_3150_out0;
assign v$RM_3531_out0 = v$_6811_out0;
assign v$RM_3532_out0 = v$_479_out0;
assign v$RM_3533_out0 = v$_3096_out0;
assign v$RM_3743_out0 = v$_7670_out0;
assign v$RM_3744_out0 = v$_8795_out0;
assign v$RM_3746_out0 = v$_10745_out0;
assign v$RM_3747_out0 = v$_13474_out0;
assign v$RM_3748_out0 = v$_8725_out0;
assign v$RM_3749_out0 = v$_3077_out0;
assign v$RM_3750_out0 = v$_3887_out0;
assign v$RM_3751_out0 = v$_3849_out0;
assign v$RM_3752_out0 = v$_2181_out0;
assign v$RM_3753_out0 = v$_1799_out0;
assign v$RM_3754_out0 = v$_3165_out0;
assign v$RM_3755_out0 = v$_6826_out0;
assign v$RM_3756_out0 = v$_494_out0;
assign v$RM_3757_out0 = v$_3111_out0;
assign v$CIN_9974_out0 = v$_2205_out0;
assign v$CIN_10198_out0 = v$_2219_out0;
assign v$RM_11654_out0 = v$_2513_out0;
assign v$RM_12118_out0 = v$_2528_out0;
assign v$RD_6207_out0 = v$CIN_9974_out0;
assign v$RD_6671_out0 = v$CIN_10198_out0;
assign v$G1_8069_out0 = ((v$RD_6214_out0 && !v$RM_11654_out0) || (!v$RD_6214_out0) && v$RM_11654_out0);
assign v$G1_8533_out0 = ((v$RD_6678_out0 && !v$RM_12118_out0) || (!v$RD_6678_out0) && v$RM_12118_out0);
assign v$RM_11642_out0 = v$RM_3519_out0;
assign v$RM_11644_out0 = v$RM_3520_out0;
assign v$RM_11648_out0 = v$RM_3522_out0;
assign v$RM_11650_out0 = v$RM_3523_out0;
assign v$RM_11652_out0 = v$RM_3524_out0;
assign v$RM_11655_out0 = v$RM_3525_out0;
assign v$RM_11657_out0 = v$RM_3526_out0;
assign v$RM_11659_out0 = v$RM_3527_out0;
assign v$RM_11661_out0 = v$RM_3528_out0;
assign v$RM_11663_out0 = v$RM_3529_out0;
assign v$RM_11665_out0 = v$RM_3530_out0;
assign v$RM_11667_out0 = v$RM_3531_out0;
assign v$RM_11669_out0 = v$RM_3532_out0;
assign v$RM_11671_out0 = v$RM_3533_out0;
assign v$RM_12106_out0 = v$RM_3743_out0;
assign v$RM_12108_out0 = v$RM_3744_out0;
assign v$RM_12112_out0 = v$RM_3746_out0;
assign v$RM_12114_out0 = v$RM_3747_out0;
assign v$RM_12116_out0 = v$RM_3748_out0;
assign v$RM_12119_out0 = v$RM_3749_out0;
assign v$RM_12121_out0 = v$RM_3750_out0;
assign v$RM_12123_out0 = v$RM_3751_out0;
assign v$RM_12125_out0 = v$RM_3752_out0;
assign v$RM_12127_out0 = v$RM_3753_out0;
assign v$RM_12129_out0 = v$RM_3754_out0;
assign v$RM_12131_out0 = v$RM_3755_out0;
assign v$RM_12133_out0 = v$RM_3756_out0;
assign v$RM_12135_out0 = v$RM_3757_out0;
assign v$G2_12605_out0 = v$RD_6214_out0 && v$RM_11654_out0;
assign v$G2_13069_out0 = v$RD_6678_out0 && v$RM_12118_out0;
assign v$CARRY_5214_out0 = v$G2_12605_out0;
assign v$CARRY_5678_out0 = v$G2_13069_out0;
assign v$G1_8057_out0 = ((v$RD_6202_out0 && !v$RM_11642_out0) || (!v$RD_6202_out0) && v$RM_11642_out0);
assign v$G1_8059_out0 = ((v$RD_6204_out0 && !v$RM_11644_out0) || (!v$RD_6204_out0) && v$RM_11644_out0);
assign v$G1_8063_out0 = ((v$RD_6208_out0 && !v$RM_11648_out0) || (!v$RD_6208_out0) && v$RM_11648_out0);
assign v$G1_8065_out0 = ((v$RD_6210_out0 && !v$RM_11650_out0) || (!v$RD_6210_out0) && v$RM_11650_out0);
assign v$G1_8067_out0 = ((v$RD_6212_out0 && !v$RM_11652_out0) || (!v$RD_6212_out0) && v$RM_11652_out0);
assign v$G1_8070_out0 = ((v$RD_6215_out0 && !v$RM_11655_out0) || (!v$RD_6215_out0) && v$RM_11655_out0);
assign v$G1_8072_out0 = ((v$RD_6217_out0 && !v$RM_11657_out0) || (!v$RD_6217_out0) && v$RM_11657_out0);
assign v$G1_8074_out0 = ((v$RD_6219_out0 && !v$RM_11659_out0) || (!v$RD_6219_out0) && v$RM_11659_out0);
assign v$G1_8076_out0 = ((v$RD_6221_out0 && !v$RM_11661_out0) || (!v$RD_6221_out0) && v$RM_11661_out0);
assign v$G1_8078_out0 = ((v$RD_6223_out0 && !v$RM_11663_out0) || (!v$RD_6223_out0) && v$RM_11663_out0);
assign v$G1_8080_out0 = ((v$RD_6225_out0 && !v$RM_11665_out0) || (!v$RD_6225_out0) && v$RM_11665_out0);
assign v$G1_8082_out0 = ((v$RD_6227_out0 && !v$RM_11667_out0) || (!v$RD_6227_out0) && v$RM_11667_out0);
assign v$G1_8084_out0 = ((v$RD_6229_out0 && !v$RM_11669_out0) || (!v$RD_6229_out0) && v$RM_11669_out0);
assign v$G1_8086_out0 = ((v$RD_6231_out0 && !v$RM_11671_out0) || (!v$RD_6231_out0) && v$RM_11671_out0);
assign v$G1_8521_out0 = ((v$RD_6666_out0 && !v$RM_12106_out0) || (!v$RD_6666_out0) && v$RM_12106_out0);
assign v$G1_8523_out0 = ((v$RD_6668_out0 && !v$RM_12108_out0) || (!v$RD_6668_out0) && v$RM_12108_out0);
assign v$G1_8527_out0 = ((v$RD_6672_out0 && !v$RM_12112_out0) || (!v$RD_6672_out0) && v$RM_12112_out0);
assign v$G1_8529_out0 = ((v$RD_6674_out0 && !v$RM_12114_out0) || (!v$RD_6674_out0) && v$RM_12114_out0);
assign v$G1_8531_out0 = ((v$RD_6676_out0 && !v$RM_12116_out0) || (!v$RD_6676_out0) && v$RM_12116_out0);
assign v$G1_8534_out0 = ((v$RD_6679_out0 && !v$RM_12119_out0) || (!v$RD_6679_out0) && v$RM_12119_out0);
assign v$G1_8536_out0 = ((v$RD_6681_out0 && !v$RM_12121_out0) || (!v$RD_6681_out0) && v$RM_12121_out0);
assign v$G1_8538_out0 = ((v$RD_6683_out0 && !v$RM_12123_out0) || (!v$RD_6683_out0) && v$RM_12123_out0);
assign v$G1_8540_out0 = ((v$RD_6685_out0 && !v$RM_12125_out0) || (!v$RD_6685_out0) && v$RM_12125_out0);
assign v$G1_8542_out0 = ((v$RD_6687_out0 && !v$RM_12127_out0) || (!v$RD_6687_out0) && v$RM_12127_out0);
assign v$G1_8544_out0 = ((v$RD_6689_out0 && !v$RM_12129_out0) || (!v$RD_6689_out0) && v$RM_12129_out0);
assign v$G1_8546_out0 = ((v$RD_6691_out0 && !v$RM_12131_out0) || (!v$RD_6691_out0) && v$RM_12131_out0);
assign v$G1_8548_out0 = ((v$RD_6693_out0 && !v$RM_12133_out0) || (!v$RD_6693_out0) && v$RM_12133_out0);
assign v$G1_8550_out0 = ((v$RD_6695_out0 && !v$RM_12135_out0) || (!v$RD_6695_out0) && v$RM_12135_out0);
assign v$S_9215_out0 = v$G1_8069_out0;
assign v$S_9679_out0 = v$G1_8533_out0;
assign v$G2_12593_out0 = v$RD_6202_out0 && v$RM_11642_out0;
assign v$G2_12595_out0 = v$RD_6204_out0 && v$RM_11644_out0;
assign v$G2_12599_out0 = v$RD_6208_out0 && v$RM_11648_out0;
assign v$G2_12601_out0 = v$RD_6210_out0 && v$RM_11650_out0;
assign v$G2_12603_out0 = v$RD_6212_out0 && v$RM_11652_out0;
assign v$G2_12606_out0 = v$RD_6215_out0 && v$RM_11655_out0;
assign v$G2_12608_out0 = v$RD_6217_out0 && v$RM_11657_out0;
assign v$G2_12610_out0 = v$RD_6219_out0 && v$RM_11659_out0;
assign v$G2_12612_out0 = v$RD_6221_out0 && v$RM_11661_out0;
assign v$G2_12614_out0 = v$RD_6223_out0 && v$RM_11663_out0;
assign v$G2_12616_out0 = v$RD_6225_out0 && v$RM_11665_out0;
assign v$G2_12618_out0 = v$RD_6227_out0 && v$RM_11667_out0;
assign v$G2_12620_out0 = v$RD_6229_out0 && v$RM_11669_out0;
assign v$G2_12622_out0 = v$RD_6231_out0 && v$RM_11671_out0;
assign v$G2_13057_out0 = v$RD_6666_out0 && v$RM_12106_out0;
assign v$G2_13059_out0 = v$RD_6668_out0 && v$RM_12108_out0;
assign v$G2_13063_out0 = v$RD_6672_out0 && v$RM_12112_out0;
assign v$G2_13065_out0 = v$RD_6674_out0 && v$RM_12114_out0;
assign v$G2_13067_out0 = v$RD_6676_out0 && v$RM_12116_out0;
assign v$G2_13070_out0 = v$RD_6679_out0 && v$RM_12119_out0;
assign v$G2_13072_out0 = v$RD_6681_out0 && v$RM_12121_out0;
assign v$G2_13074_out0 = v$RD_6683_out0 && v$RM_12123_out0;
assign v$G2_13076_out0 = v$RD_6685_out0 && v$RM_12125_out0;
assign v$G2_13078_out0 = v$RD_6687_out0 && v$RM_12127_out0;
assign v$G2_13080_out0 = v$RD_6689_out0 && v$RM_12129_out0;
assign v$G2_13082_out0 = v$RD_6691_out0 && v$RM_12131_out0;
assign v$G2_13084_out0 = v$RD_6693_out0 && v$RM_12133_out0;
assign v$G2_13086_out0 = v$RD_6695_out0 && v$RM_12135_out0;
assign v$S_4676_out0 = v$S_9215_out0;
assign v$S_4691_out0 = v$S_9679_out0;
assign v$CARRY_5202_out0 = v$G2_12593_out0;
assign v$CARRY_5204_out0 = v$G2_12595_out0;
assign v$CARRY_5208_out0 = v$G2_12599_out0;
assign v$CARRY_5210_out0 = v$G2_12601_out0;
assign v$CARRY_5212_out0 = v$G2_12603_out0;
assign v$CARRY_5215_out0 = v$G2_12606_out0;
assign v$CARRY_5217_out0 = v$G2_12608_out0;
assign v$CARRY_5219_out0 = v$G2_12610_out0;
assign v$CARRY_5221_out0 = v$G2_12612_out0;
assign v$CARRY_5223_out0 = v$G2_12614_out0;
assign v$CARRY_5225_out0 = v$G2_12616_out0;
assign v$CARRY_5227_out0 = v$G2_12618_out0;
assign v$CARRY_5229_out0 = v$G2_12620_out0;
assign v$CARRY_5231_out0 = v$G2_12622_out0;
assign v$CARRY_5666_out0 = v$G2_13057_out0;
assign v$CARRY_5668_out0 = v$G2_13059_out0;
assign v$CARRY_5672_out0 = v$G2_13063_out0;
assign v$CARRY_5674_out0 = v$G2_13065_out0;
assign v$CARRY_5676_out0 = v$G2_13067_out0;
assign v$CARRY_5679_out0 = v$G2_13070_out0;
assign v$CARRY_5681_out0 = v$G2_13072_out0;
assign v$CARRY_5683_out0 = v$G2_13074_out0;
assign v$CARRY_5685_out0 = v$G2_13076_out0;
assign v$CARRY_5687_out0 = v$G2_13078_out0;
assign v$CARRY_5689_out0 = v$G2_13080_out0;
assign v$CARRY_5691_out0 = v$G2_13082_out0;
assign v$CARRY_5693_out0 = v$G2_13084_out0;
assign v$CARRY_5695_out0 = v$G2_13086_out0;
assign v$S_9203_out0 = v$G1_8057_out0;
assign v$S_9205_out0 = v$G1_8059_out0;
assign v$S_9209_out0 = v$G1_8063_out0;
assign v$S_9211_out0 = v$G1_8065_out0;
assign v$S_9213_out0 = v$G1_8067_out0;
assign v$S_9216_out0 = v$G1_8070_out0;
assign v$S_9218_out0 = v$G1_8072_out0;
assign v$S_9220_out0 = v$G1_8074_out0;
assign v$S_9222_out0 = v$G1_8076_out0;
assign v$S_9224_out0 = v$G1_8078_out0;
assign v$S_9226_out0 = v$G1_8080_out0;
assign v$S_9228_out0 = v$G1_8082_out0;
assign v$S_9230_out0 = v$G1_8084_out0;
assign v$S_9232_out0 = v$G1_8086_out0;
assign v$S_9667_out0 = v$G1_8521_out0;
assign v$S_9669_out0 = v$G1_8523_out0;
assign v$S_9673_out0 = v$G1_8527_out0;
assign v$S_9675_out0 = v$G1_8529_out0;
assign v$S_9677_out0 = v$G1_8531_out0;
assign v$S_9680_out0 = v$G1_8534_out0;
assign v$S_9682_out0 = v$G1_8536_out0;
assign v$S_9684_out0 = v$G1_8538_out0;
assign v$S_9686_out0 = v$G1_8540_out0;
assign v$S_9688_out0 = v$G1_8542_out0;
assign v$S_9690_out0 = v$G1_8544_out0;
assign v$S_9692_out0 = v$G1_8546_out0;
assign v$S_9694_out0 = v$G1_8548_out0;
assign v$S_9696_out0 = v$G1_8550_out0;
assign v$CIN_9980_out0 = v$CARRY_5214_out0;
assign v$CIN_10204_out0 = v$CARRY_5678_out0;
assign v$_636_out0 = { v$_681_out0,v$S_4676_out0 };
assign v$_637_out0 = { v$_682_out0,v$S_4691_out0 };
assign v$RD_6220_out0 = v$CIN_9980_out0;
assign v$RD_6684_out0 = v$CIN_10204_out0;
assign v$RM_11643_out0 = v$S_9203_out0;
assign v$RM_11645_out0 = v$S_9205_out0;
assign v$RM_11649_out0 = v$S_9209_out0;
assign v$RM_11651_out0 = v$S_9211_out0;
assign v$RM_11653_out0 = v$S_9213_out0;
assign v$RM_11656_out0 = v$S_9216_out0;
assign v$RM_11658_out0 = v$S_9218_out0;
assign v$RM_11660_out0 = v$S_9220_out0;
assign v$RM_11662_out0 = v$S_9222_out0;
assign v$RM_11664_out0 = v$S_9224_out0;
assign v$RM_11666_out0 = v$S_9226_out0;
assign v$RM_11668_out0 = v$S_9228_out0;
assign v$RM_11670_out0 = v$S_9230_out0;
assign v$RM_11672_out0 = v$S_9232_out0;
assign v$RM_12107_out0 = v$S_9667_out0;
assign v$RM_12109_out0 = v$S_9669_out0;
assign v$RM_12113_out0 = v$S_9673_out0;
assign v$RM_12115_out0 = v$S_9675_out0;
assign v$RM_12117_out0 = v$S_9677_out0;
assign v$RM_12120_out0 = v$S_9680_out0;
assign v$RM_12122_out0 = v$S_9682_out0;
assign v$RM_12124_out0 = v$S_9684_out0;
assign v$RM_12126_out0 = v$S_9686_out0;
assign v$RM_12128_out0 = v$S_9688_out0;
assign v$RM_12130_out0 = v$S_9690_out0;
assign v$RM_12132_out0 = v$S_9692_out0;
assign v$RM_12134_out0 = v$S_9694_out0;
assign v$RM_12136_out0 = v$S_9696_out0;
assign v$G1_8075_out0 = ((v$RD_6220_out0 && !v$RM_11660_out0) || (!v$RD_6220_out0) && v$RM_11660_out0);
assign v$G1_8539_out0 = ((v$RD_6684_out0 && !v$RM_12124_out0) || (!v$RD_6684_out0) && v$RM_12124_out0);
assign v$G2_12611_out0 = v$RD_6220_out0 && v$RM_11660_out0;
assign v$G2_13075_out0 = v$RD_6684_out0 && v$RM_12124_out0;
assign v$CARRY_5220_out0 = v$G2_12611_out0;
assign v$CARRY_5684_out0 = v$G2_13075_out0;
assign v$S_9221_out0 = v$G1_8075_out0;
assign v$S_9685_out0 = v$G1_8539_out0;
assign v$S_1391_out0 = v$S_9221_out0;
assign v$S_1615_out0 = v$S_9685_out0;
assign v$G1_4167_out0 = v$CARRY_5220_out0 || v$CARRY_5219_out0;
assign v$G1_4391_out0 = v$CARRY_5684_out0 || v$CARRY_5683_out0;
assign v$COUT_859_out0 = v$G1_4167_out0;
assign v$COUT_1083_out0 = v$G1_4391_out0;
assign v$CIN_9986_out0 = v$COUT_859_out0;
assign v$CIN_10210_out0 = v$COUT_1083_out0;
assign v$RD_6232_out0 = v$CIN_9986_out0;
assign v$RD_6696_out0 = v$CIN_10210_out0;
assign v$G1_8087_out0 = ((v$RD_6232_out0 && !v$RM_11672_out0) || (!v$RD_6232_out0) && v$RM_11672_out0);
assign v$G1_8551_out0 = ((v$RD_6696_out0 && !v$RM_12136_out0) || (!v$RD_6696_out0) && v$RM_12136_out0);
assign v$G2_12623_out0 = v$RD_6232_out0 && v$RM_11672_out0;
assign v$G2_13087_out0 = v$RD_6696_out0 && v$RM_12136_out0;
assign v$CARRY_5232_out0 = v$G2_12623_out0;
assign v$CARRY_5696_out0 = v$G2_13087_out0;
assign v$S_9233_out0 = v$G1_8087_out0;
assign v$S_9697_out0 = v$G1_8551_out0;
assign v$S_1397_out0 = v$S_9233_out0;
assign v$S_1621_out0 = v$S_9697_out0;
assign v$G1_4173_out0 = v$CARRY_5232_out0 || v$CARRY_5231_out0;
assign v$G1_4397_out0 = v$CARRY_5696_out0 || v$CARRY_5695_out0;
assign v$COUT_865_out0 = v$G1_4173_out0;
assign v$COUT_1089_out0 = v$G1_4397_out0;
assign v$_4793_out0 = { v$S_1391_out0,v$S_1397_out0 };
assign v$_4808_out0 = { v$S_1615_out0,v$S_1621_out0 };
assign v$CIN_9981_out0 = v$COUT_865_out0;
assign v$CIN_10205_out0 = v$COUT_1089_out0;
assign v$RD_6222_out0 = v$CIN_9981_out0;
assign v$RD_6686_out0 = v$CIN_10205_out0;
assign v$G1_8077_out0 = ((v$RD_6222_out0 && !v$RM_11662_out0) || (!v$RD_6222_out0) && v$RM_11662_out0);
assign v$G1_8541_out0 = ((v$RD_6686_out0 && !v$RM_12126_out0) || (!v$RD_6686_out0) && v$RM_12126_out0);
assign v$G2_12613_out0 = v$RD_6222_out0 && v$RM_11662_out0;
assign v$G2_13077_out0 = v$RD_6686_out0 && v$RM_12126_out0;
assign v$CARRY_5222_out0 = v$G2_12613_out0;
assign v$CARRY_5686_out0 = v$G2_13077_out0;
assign v$S_9223_out0 = v$G1_8077_out0;
assign v$S_9687_out0 = v$G1_8541_out0;
assign v$S_1392_out0 = v$S_9223_out0;
assign v$S_1616_out0 = v$S_9687_out0;
assign v$G1_4168_out0 = v$CARRY_5222_out0 || v$CARRY_5221_out0;
assign v$G1_4392_out0 = v$CARRY_5686_out0 || v$CARRY_5685_out0;
assign v$COUT_860_out0 = v$G1_4168_out0;
assign v$COUT_1084_out0 = v$G1_4392_out0;
assign v$_2563_out0 = { v$_4793_out0,v$S_1392_out0 };
assign v$_2578_out0 = { v$_4808_out0,v$S_1616_out0 };
assign v$CIN_9976_out0 = v$COUT_860_out0;
assign v$CIN_10200_out0 = v$COUT_1084_out0;
assign v$RD_6211_out0 = v$CIN_9976_out0;
assign v$RD_6675_out0 = v$CIN_10200_out0;
assign v$G1_8066_out0 = ((v$RD_6211_out0 && !v$RM_11651_out0) || (!v$RD_6211_out0) && v$RM_11651_out0);
assign v$G1_8530_out0 = ((v$RD_6675_out0 && !v$RM_12115_out0) || (!v$RD_6675_out0) && v$RM_12115_out0);
assign v$G2_12602_out0 = v$RD_6211_out0 && v$RM_11651_out0;
assign v$G2_13066_out0 = v$RD_6675_out0 && v$RM_12115_out0;
assign v$CARRY_5211_out0 = v$G2_12602_out0;
assign v$CARRY_5675_out0 = v$G2_13066_out0;
assign v$S_9212_out0 = v$G1_8066_out0;
assign v$S_9676_out0 = v$G1_8530_out0;
assign v$S_1387_out0 = v$S_9212_out0;
assign v$S_1611_out0 = v$S_9676_out0;
assign v$G1_4163_out0 = v$CARRY_5211_out0 || v$CARRY_5210_out0;
assign v$G1_4387_out0 = v$CARRY_5675_out0 || v$CARRY_5674_out0;
assign v$COUT_855_out0 = v$G1_4163_out0;
assign v$COUT_1079_out0 = v$G1_4387_out0;
assign v$_7043_out0 = { v$_2563_out0,v$S_1387_out0 };
assign v$_7058_out0 = { v$_2578_out0,v$S_1611_out0 };
assign v$CIN_9975_out0 = v$COUT_855_out0;
assign v$CIN_10199_out0 = v$COUT_1079_out0;
assign v$RD_6209_out0 = v$CIN_9975_out0;
assign v$RD_6673_out0 = v$CIN_10199_out0;
assign v$G1_8064_out0 = ((v$RD_6209_out0 && !v$RM_11649_out0) || (!v$RD_6209_out0) && v$RM_11649_out0);
assign v$G1_8528_out0 = ((v$RD_6673_out0 && !v$RM_12113_out0) || (!v$RD_6673_out0) && v$RM_12113_out0);
assign v$G2_12600_out0 = v$RD_6209_out0 && v$RM_11649_out0;
assign v$G2_13064_out0 = v$RD_6673_out0 && v$RM_12113_out0;
assign v$CARRY_5209_out0 = v$G2_12600_out0;
assign v$CARRY_5673_out0 = v$G2_13064_out0;
assign v$S_9210_out0 = v$G1_8064_out0;
assign v$S_9674_out0 = v$G1_8528_out0;
assign v$S_1386_out0 = v$S_9210_out0;
assign v$S_1610_out0 = v$S_9674_out0;
assign v$G1_4162_out0 = v$CARRY_5209_out0 || v$CARRY_5208_out0;
assign v$G1_4386_out0 = v$CARRY_5673_out0 || v$CARRY_5672_out0;
assign v$COUT_854_out0 = v$G1_4162_out0;
assign v$COUT_1078_out0 = v$G1_4386_out0;
assign v$_13529_out0 = { v$_7043_out0,v$S_1386_out0 };
assign v$_13544_out0 = { v$_7058_out0,v$S_1610_out0 };
assign v$CIN_9982_out0 = v$COUT_854_out0;
assign v$CIN_10206_out0 = v$COUT_1078_out0;
assign v$RD_6224_out0 = v$CIN_9982_out0;
assign v$RD_6688_out0 = v$CIN_10206_out0;
assign v$G1_8079_out0 = ((v$RD_6224_out0 && !v$RM_11664_out0) || (!v$RD_6224_out0) && v$RM_11664_out0);
assign v$G1_8543_out0 = ((v$RD_6688_out0 && !v$RM_12128_out0) || (!v$RD_6688_out0) && v$RM_12128_out0);
assign v$G2_12615_out0 = v$RD_6224_out0 && v$RM_11664_out0;
assign v$G2_13079_out0 = v$RD_6688_out0 && v$RM_12128_out0;
assign v$CARRY_5224_out0 = v$G2_12615_out0;
assign v$CARRY_5688_out0 = v$G2_13079_out0;
assign v$S_9225_out0 = v$G1_8079_out0;
assign v$S_9689_out0 = v$G1_8543_out0;
assign v$S_1393_out0 = v$S_9225_out0;
assign v$S_1617_out0 = v$S_9689_out0;
assign v$G1_4169_out0 = v$CARRY_5224_out0 || v$CARRY_5223_out0;
assign v$G1_4393_out0 = v$CARRY_5688_out0 || v$CARRY_5687_out0;
assign v$COUT_861_out0 = v$G1_4169_out0;
assign v$COUT_1085_out0 = v$G1_4393_out0;
assign v$_3322_out0 = { v$_13529_out0,v$S_1393_out0 };
assign v$_3337_out0 = { v$_13544_out0,v$S_1617_out0 };
assign v$CIN_9983_out0 = v$COUT_861_out0;
assign v$CIN_10207_out0 = v$COUT_1085_out0;
assign v$RD_6226_out0 = v$CIN_9983_out0;
assign v$RD_6690_out0 = v$CIN_10207_out0;
assign v$G1_8081_out0 = ((v$RD_6226_out0 && !v$RM_11666_out0) || (!v$RD_6226_out0) && v$RM_11666_out0);
assign v$G1_8545_out0 = ((v$RD_6690_out0 && !v$RM_12130_out0) || (!v$RD_6690_out0) && v$RM_12130_out0);
assign v$G2_12617_out0 = v$RD_6226_out0 && v$RM_11666_out0;
assign v$G2_13081_out0 = v$RD_6690_out0 && v$RM_12130_out0;
assign v$CARRY_5226_out0 = v$G2_12617_out0;
assign v$CARRY_5690_out0 = v$G2_13081_out0;
assign v$S_9227_out0 = v$G1_8081_out0;
assign v$S_9691_out0 = v$G1_8545_out0;
assign v$S_1394_out0 = v$S_9227_out0;
assign v$S_1618_out0 = v$S_9691_out0;
assign v$G1_4170_out0 = v$CARRY_5226_out0 || v$CARRY_5225_out0;
assign v$G1_4394_out0 = v$CARRY_5690_out0 || v$CARRY_5689_out0;
assign v$COUT_862_out0 = v$G1_4170_out0;
assign v$COUT_1086_out0 = v$G1_4394_out0;
assign v$_7158_out0 = { v$_3322_out0,v$S_1394_out0 };
assign v$_7173_out0 = { v$_3337_out0,v$S_1618_out0 };
assign v$CIN_9985_out0 = v$COUT_862_out0;
assign v$CIN_10209_out0 = v$COUT_1086_out0;
assign v$RD_6230_out0 = v$CIN_9985_out0;
assign v$RD_6694_out0 = v$CIN_10209_out0;
assign v$G1_8085_out0 = ((v$RD_6230_out0 && !v$RM_11670_out0) || (!v$RD_6230_out0) && v$RM_11670_out0);
assign v$G1_8549_out0 = ((v$RD_6694_out0 && !v$RM_12134_out0) || (!v$RD_6694_out0) && v$RM_12134_out0);
assign v$G2_12621_out0 = v$RD_6230_out0 && v$RM_11670_out0;
assign v$G2_13085_out0 = v$RD_6694_out0 && v$RM_12134_out0;
assign v$CARRY_5230_out0 = v$G2_12621_out0;
assign v$CARRY_5694_out0 = v$G2_13085_out0;
assign v$S_9231_out0 = v$G1_8085_out0;
assign v$S_9695_out0 = v$G1_8549_out0;
assign v$S_1396_out0 = v$S_9231_out0;
assign v$S_1620_out0 = v$S_9695_out0;
assign v$G1_4172_out0 = v$CARRY_5230_out0 || v$CARRY_5229_out0;
assign v$G1_4396_out0 = v$CARRY_5694_out0 || v$CARRY_5693_out0;
assign v$COUT_864_out0 = v$G1_4172_out0;
assign v$COUT_1088_out0 = v$G1_4396_out0;
assign v$_4760_out0 = { v$_7158_out0,v$S_1396_out0 };
assign v$_4775_out0 = { v$_7173_out0,v$S_1620_out0 };
assign v$CIN_9978_out0 = v$COUT_864_out0;
assign v$CIN_10202_out0 = v$COUT_1088_out0;
assign v$RD_6216_out0 = v$CIN_9978_out0;
assign v$RD_6680_out0 = v$CIN_10202_out0;
assign v$G1_8071_out0 = ((v$RD_6216_out0 && !v$RM_11656_out0) || (!v$RD_6216_out0) && v$RM_11656_out0);
assign v$G1_8535_out0 = ((v$RD_6680_out0 && !v$RM_12120_out0) || (!v$RD_6680_out0) && v$RM_12120_out0);
assign v$G2_12607_out0 = v$RD_6216_out0 && v$RM_11656_out0;
assign v$G2_13071_out0 = v$RD_6680_out0 && v$RM_12120_out0;
assign v$CARRY_5216_out0 = v$G2_12607_out0;
assign v$CARRY_5680_out0 = v$G2_13071_out0;
assign v$S_9217_out0 = v$G1_8071_out0;
assign v$S_9681_out0 = v$G1_8535_out0;
assign v$S_1389_out0 = v$S_9217_out0;
assign v$S_1613_out0 = v$S_9681_out0;
assign v$G1_4165_out0 = v$CARRY_5216_out0 || v$CARRY_5215_out0;
assign v$G1_4389_out0 = v$CARRY_5680_out0 || v$CARRY_5679_out0;
assign v$COUT_857_out0 = v$G1_4165_out0;
assign v$COUT_1081_out0 = v$G1_4389_out0;
assign v$_6937_out0 = { v$_4760_out0,v$S_1389_out0 };
assign v$_6952_out0 = { v$_4775_out0,v$S_1613_out0 };
assign v$CIN_9979_out0 = v$COUT_857_out0;
assign v$CIN_10203_out0 = v$COUT_1081_out0;
assign v$RD_6218_out0 = v$CIN_9979_out0;
assign v$RD_6682_out0 = v$CIN_10203_out0;
assign v$G1_8073_out0 = ((v$RD_6218_out0 && !v$RM_11658_out0) || (!v$RD_6218_out0) && v$RM_11658_out0);
assign v$G1_8537_out0 = ((v$RD_6682_out0 && !v$RM_12122_out0) || (!v$RD_6682_out0) && v$RM_12122_out0);
assign v$G2_12609_out0 = v$RD_6218_out0 && v$RM_11658_out0;
assign v$G2_13073_out0 = v$RD_6682_out0 && v$RM_12122_out0;
assign v$CARRY_5218_out0 = v$G2_12609_out0;
assign v$CARRY_5682_out0 = v$G2_13073_out0;
assign v$S_9219_out0 = v$G1_8073_out0;
assign v$S_9683_out0 = v$G1_8537_out0;
assign v$S_1390_out0 = v$S_9219_out0;
assign v$S_1614_out0 = v$S_9683_out0;
assign v$G1_4166_out0 = v$CARRY_5218_out0 || v$CARRY_5217_out0;
assign v$G1_4390_out0 = v$CARRY_5682_out0 || v$CARRY_5681_out0;
assign v$COUT_858_out0 = v$G1_4166_out0;
assign v$COUT_1082_out0 = v$G1_4390_out0;
assign v$_5813_out0 = { v$_6937_out0,v$S_1390_out0 };
assign v$_5828_out0 = { v$_6952_out0,v$S_1614_out0 };
assign v$CIN_9984_out0 = v$COUT_858_out0;
assign v$CIN_10208_out0 = v$COUT_1082_out0;
assign v$RD_6228_out0 = v$CIN_9984_out0;
assign v$RD_6692_out0 = v$CIN_10208_out0;
assign v$G1_8083_out0 = ((v$RD_6228_out0 && !v$RM_11668_out0) || (!v$RD_6228_out0) && v$RM_11668_out0);
assign v$G1_8547_out0 = ((v$RD_6692_out0 && !v$RM_12132_out0) || (!v$RD_6692_out0) && v$RM_12132_out0);
assign v$G2_12619_out0 = v$RD_6228_out0 && v$RM_11668_out0;
assign v$G2_13083_out0 = v$RD_6692_out0 && v$RM_12132_out0;
assign v$CARRY_5228_out0 = v$G2_12619_out0;
assign v$CARRY_5692_out0 = v$G2_13083_out0;
assign v$S_9229_out0 = v$G1_8083_out0;
assign v$S_9693_out0 = v$G1_8547_out0;
assign v$S_1395_out0 = v$S_9229_out0;
assign v$S_1619_out0 = v$S_9693_out0;
assign v$G1_4171_out0 = v$CARRY_5228_out0 || v$CARRY_5227_out0;
assign v$G1_4395_out0 = v$CARRY_5692_out0 || v$CARRY_5691_out0;
assign v$COUT_863_out0 = v$G1_4171_out0;
assign v$COUT_1087_out0 = v$G1_4395_out0;
assign v$_2037_out0 = { v$_5813_out0,v$S_1395_out0 };
assign v$_2052_out0 = { v$_5828_out0,v$S_1619_out0 };
assign v$CIN_9972_out0 = v$COUT_863_out0;
assign v$CIN_10196_out0 = v$COUT_1087_out0;
assign v$RD_6203_out0 = v$CIN_9972_out0;
assign v$RD_6667_out0 = v$CIN_10196_out0;
assign v$G1_8058_out0 = ((v$RD_6203_out0 && !v$RM_11643_out0) || (!v$RD_6203_out0) && v$RM_11643_out0);
assign v$G1_8522_out0 = ((v$RD_6667_out0 && !v$RM_12107_out0) || (!v$RD_6667_out0) && v$RM_12107_out0);
assign v$G2_12594_out0 = v$RD_6203_out0 && v$RM_11643_out0;
assign v$G2_13058_out0 = v$RD_6667_out0 && v$RM_12107_out0;
assign v$CARRY_5203_out0 = v$G2_12594_out0;
assign v$CARRY_5667_out0 = v$G2_13058_out0;
assign v$S_9204_out0 = v$G1_8058_out0;
assign v$S_9668_out0 = v$G1_8522_out0;
assign v$S_1383_out0 = v$S_9204_out0;
assign v$S_1607_out0 = v$S_9668_out0;
assign v$G1_4159_out0 = v$CARRY_5203_out0 || v$CARRY_5202_out0;
assign v$G1_4383_out0 = v$CARRY_5667_out0 || v$CARRY_5666_out0;
assign v$COUT_851_out0 = v$G1_4159_out0;
assign v$COUT_1075_out0 = v$G1_4383_out0;
assign v$_2804_out0 = { v$_2037_out0,v$S_1383_out0 };
assign v$_2819_out0 = { v$_2052_out0,v$S_1607_out0 };
assign v$CIN_9977_out0 = v$COUT_851_out0;
assign v$CIN_10201_out0 = v$COUT_1075_out0;
assign v$RD_6213_out0 = v$CIN_9977_out0;
assign v$RD_6677_out0 = v$CIN_10201_out0;
assign v$G1_8068_out0 = ((v$RD_6213_out0 && !v$RM_11653_out0) || (!v$RD_6213_out0) && v$RM_11653_out0);
assign v$G1_8532_out0 = ((v$RD_6677_out0 && !v$RM_12117_out0) || (!v$RD_6677_out0) && v$RM_12117_out0);
assign v$G2_12604_out0 = v$RD_6213_out0 && v$RM_11653_out0;
assign v$G2_13068_out0 = v$RD_6677_out0 && v$RM_12117_out0;
assign v$CARRY_5213_out0 = v$G2_12604_out0;
assign v$CARRY_5677_out0 = v$G2_13068_out0;
assign v$S_9214_out0 = v$G1_8068_out0;
assign v$S_9678_out0 = v$G1_8532_out0;
assign v$S_1388_out0 = v$S_9214_out0;
assign v$S_1612_out0 = v$S_9678_out0;
assign v$G1_4164_out0 = v$CARRY_5213_out0 || v$CARRY_5212_out0;
assign v$G1_4388_out0 = v$CARRY_5677_out0 || v$CARRY_5676_out0;
assign v$COUT_856_out0 = v$G1_4164_out0;
assign v$COUT_1080_out0 = v$G1_4388_out0;
assign v$_1836_out0 = { v$_2804_out0,v$S_1388_out0 };
assign v$_1851_out0 = { v$_2819_out0,v$S_1612_out0 };
assign v$CIN_9973_out0 = v$COUT_856_out0;
assign v$CIN_10197_out0 = v$COUT_1080_out0;
assign v$RD_6205_out0 = v$CIN_9973_out0;
assign v$RD_6669_out0 = v$CIN_10197_out0;
assign v$G1_8060_out0 = ((v$RD_6205_out0 && !v$RM_11645_out0) || (!v$RD_6205_out0) && v$RM_11645_out0);
assign v$G1_8524_out0 = ((v$RD_6669_out0 && !v$RM_12109_out0) || (!v$RD_6669_out0) && v$RM_12109_out0);
assign v$G2_12596_out0 = v$RD_6205_out0 && v$RM_11645_out0;
assign v$G2_13060_out0 = v$RD_6669_out0 && v$RM_12109_out0;
assign v$CARRY_5205_out0 = v$G2_12596_out0;
assign v$CARRY_5669_out0 = v$G2_13060_out0;
assign v$S_9206_out0 = v$G1_8060_out0;
assign v$S_9670_out0 = v$G1_8524_out0;
assign v$S_1384_out0 = v$S_9206_out0;
assign v$S_1608_out0 = v$S_9670_out0;
assign v$G1_4160_out0 = v$CARRY_5205_out0 || v$CARRY_5204_out0;
assign v$G1_4384_out0 = v$CARRY_5669_out0 || v$CARRY_5668_out0;
assign v$COUT_852_out0 = v$G1_4160_out0;
assign v$COUT_1076_out0 = v$G1_4384_out0;
assign v$_4560_out0 = { v$_1836_out0,v$S_1384_out0 };
assign v$_4575_out0 = { v$_1851_out0,v$S_1608_out0 };
assign v$RM_3521_out0 = v$COUT_852_out0;
assign v$RM_3745_out0 = v$COUT_1076_out0;
assign v$RM_11646_out0 = v$RM_3521_out0;
assign v$RM_12110_out0 = v$RM_3745_out0;
assign v$G1_8061_out0 = ((v$RD_6206_out0 && !v$RM_11646_out0) || (!v$RD_6206_out0) && v$RM_11646_out0);
assign v$G1_8525_out0 = ((v$RD_6670_out0 && !v$RM_12110_out0) || (!v$RD_6670_out0) && v$RM_12110_out0);
assign v$G2_12597_out0 = v$RD_6206_out0 && v$RM_11646_out0;
assign v$G2_13061_out0 = v$RD_6670_out0 && v$RM_12110_out0;
assign v$CARRY_5206_out0 = v$G2_12597_out0;
assign v$CARRY_5670_out0 = v$G2_13061_out0;
assign v$S_9207_out0 = v$G1_8061_out0;
assign v$S_9671_out0 = v$G1_8525_out0;
assign v$RM_11647_out0 = v$S_9207_out0;
assign v$RM_12111_out0 = v$S_9671_out0;
assign v$G1_8062_out0 = ((v$RD_6207_out0 && !v$RM_11647_out0) || (!v$RD_6207_out0) && v$RM_11647_out0);
assign v$G1_8526_out0 = ((v$RD_6671_out0 && !v$RM_12111_out0) || (!v$RD_6671_out0) && v$RM_12111_out0);
assign v$G2_12598_out0 = v$RD_6207_out0 && v$RM_11647_out0;
assign v$G2_13062_out0 = v$RD_6671_out0 && v$RM_12111_out0;
assign v$CARRY_5207_out0 = v$G2_12598_out0;
assign v$CARRY_5671_out0 = v$G2_13062_out0;
assign v$S_9208_out0 = v$G1_8062_out0;
assign v$S_9672_out0 = v$G1_8526_out0;
assign v$S_1385_out0 = v$S_9208_out0;
assign v$S_1609_out0 = v$S_9672_out0;
assign v$G1_4161_out0 = v$CARRY_5207_out0 || v$CARRY_5206_out0;
assign v$G1_4385_out0 = v$CARRY_5671_out0 || v$CARRY_5670_out0;
assign v$COUT_853_out0 = v$G1_4161_out0;
assign v$COUT_1077_out0 = v$G1_4385_out0;
assign v$_10662_out0 = { v$_4560_out0,v$S_1385_out0 };
assign v$_10677_out0 = { v$_4575_out0,v$S_1609_out0 };
assign v$_10957_out0 = { v$_10662_out0,v$COUT_853_out0 };
assign v$_10972_out0 = { v$_10677_out0,v$COUT_1077_out0 };
assign v$COUT_10927_out0 = v$_10957_out0;
assign v$COUT_10942_out0 = v$_10972_out0;
assign v$CIN_2364_out0 = v$COUT_10927_out0;
assign v$CIN_2379_out0 = v$COUT_10942_out0;
assign v$_477_out0 = v$CIN_2364_out0[8:8];
assign v$_492_out0 = v$CIN_2379_out0[8:8];
assign v$_1782_out0 = v$CIN_2364_out0[6:6];
assign v$_1797_out0 = v$CIN_2379_out0[6:6];
assign v$_2164_out0 = v$CIN_2364_out0[3:3];
assign v$_2179_out0 = v$CIN_2379_out0[3:3];
assign v$_2203_out0 = v$CIN_2364_out0[15:15];
assign v$_2217_out0 = v$CIN_2379_out0[15:15];
assign v$_2511_out0 = v$CIN_2364_out0[0:0];
assign v$_2526_out0 = v$CIN_2379_out0[0:0];
assign v$_3060_out0 = v$CIN_2364_out0[9:9];
assign v$_3075_out0 = v$CIN_2379_out0[9:9];
assign v$_3094_out0 = v$CIN_2364_out0[2:2];
assign v$_3109_out0 = v$CIN_2379_out0[2:2];
assign v$_3148_out0 = v$CIN_2364_out0[7:7];
assign v$_3163_out0 = v$CIN_2379_out0[7:7];
assign v$_3832_out0 = v$CIN_2364_out0[1:1];
assign v$_3847_out0 = v$CIN_2379_out0[1:1];
assign v$_3870_out0 = v$CIN_2364_out0[10:10];
assign v$_3885_out0 = v$CIN_2379_out0[10:10];
assign v$_6809_out0 = v$CIN_2364_out0[11:11];
assign v$_6824_out0 = v$CIN_2379_out0[11:11];
assign v$_7653_out0 = v$CIN_2364_out0[12:12];
assign v$_7668_out0 = v$CIN_2379_out0[12:12];
assign v$_8708_out0 = v$CIN_2364_out0[13:13];
assign v$_8723_out0 = v$CIN_2379_out0[13:13];
assign v$_8778_out0 = v$CIN_2364_out0[14:14];
assign v$_8793_out0 = v$CIN_2379_out0[14:14];
assign v$_10728_out0 = v$CIN_2364_out0[5:5];
assign v$_10743_out0 = v$CIN_2379_out0[5:5];
assign v$_13457_out0 = v$CIN_2364_out0[4:4];
assign v$_13472_out0 = v$CIN_2379_out0[4:4];
assign v$RM_3489_out0 = v$_7653_out0;
assign v$RM_3490_out0 = v$_8778_out0;
assign v$RM_3492_out0 = v$_10728_out0;
assign v$RM_3493_out0 = v$_13457_out0;
assign v$RM_3494_out0 = v$_8708_out0;
assign v$RM_3495_out0 = v$_3060_out0;
assign v$RM_3496_out0 = v$_3870_out0;
assign v$RM_3497_out0 = v$_3832_out0;
assign v$RM_3498_out0 = v$_2164_out0;
assign v$RM_3499_out0 = v$_1782_out0;
assign v$RM_3500_out0 = v$_3148_out0;
assign v$RM_3501_out0 = v$_6809_out0;
assign v$RM_3502_out0 = v$_477_out0;
assign v$RM_3503_out0 = v$_3094_out0;
assign v$RM_3713_out0 = v$_7668_out0;
assign v$RM_3714_out0 = v$_8793_out0;
assign v$RM_3716_out0 = v$_10743_out0;
assign v$RM_3717_out0 = v$_13472_out0;
assign v$RM_3718_out0 = v$_8723_out0;
assign v$RM_3719_out0 = v$_3075_out0;
assign v$RM_3720_out0 = v$_3885_out0;
assign v$RM_3721_out0 = v$_3847_out0;
assign v$RM_3722_out0 = v$_2179_out0;
assign v$RM_3723_out0 = v$_1797_out0;
assign v$RM_3724_out0 = v$_3163_out0;
assign v$RM_3725_out0 = v$_6824_out0;
assign v$RM_3726_out0 = v$_492_out0;
assign v$RM_3727_out0 = v$_3109_out0;
assign v$CIN_9944_out0 = v$_2203_out0;
assign v$CIN_10168_out0 = v$_2217_out0;
assign v$RM_11592_out0 = v$_2511_out0;
assign v$RM_12056_out0 = v$_2526_out0;
assign v$RD_6145_out0 = v$CIN_9944_out0;
assign v$RD_6609_out0 = v$CIN_10168_out0;
assign v$G1_8007_out0 = ((v$RD_6152_out0 && !v$RM_11592_out0) || (!v$RD_6152_out0) && v$RM_11592_out0);
assign v$G1_8471_out0 = ((v$RD_6616_out0 && !v$RM_12056_out0) || (!v$RD_6616_out0) && v$RM_12056_out0);
assign v$RM_11580_out0 = v$RM_3489_out0;
assign v$RM_11582_out0 = v$RM_3490_out0;
assign v$RM_11586_out0 = v$RM_3492_out0;
assign v$RM_11588_out0 = v$RM_3493_out0;
assign v$RM_11590_out0 = v$RM_3494_out0;
assign v$RM_11593_out0 = v$RM_3495_out0;
assign v$RM_11595_out0 = v$RM_3496_out0;
assign v$RM_11597_out0 = v$RM_3497_out0;
assign v$RM_11599_out0 = v$RM_3498_out0;
assign v$RM_11601_out0 = v$RM_3499_out0;
assign v$RM_11603_out0 = v$RM_3500_out0;
assign v$RM_11605_out0 = v$RM_3501_out0;
assign v$RM_11607_out0 = v$RM_3502_out0;
assign v$RM_11609_out0 = v$RM_3503_out0;
assign v$RM_12044_out0 = v$RM_3713_out0;
assign v$RM_12046_out0 = v$RM_3714_out0;
assign v$RM_12050_out0 = v$RM_3716_out0;
assign v$RM_12052_out0 = v$RM_3717_out0;
assign v$RM_12054_out0 = v$RM_3718_out0;
assign v$RM_12057_out0 = v$RM_3719_out0;
assign v$RM_12059_out0 = v$RM_3720_out0;
assign v$RM_12061_out0 = v$RM_3721_out0;
assign v$RM_12063_out0 = v$RM_3722_out0;
assign v$RM_12065_out0 = v$RM_3723_out0;
assign v$RM_12067_out0 = v$RM_3724_out0;
assign v$RM_12069_out0 = v$RM_3725_out0;
assign v$RM_12071_out0 = v$RM_3726_out0;
assign v$RM_12073_out0 = v$RM_3727_out0;
assign v$G2_12543_out0 = v$RD_6152_out0 && v$RM_11592_out0;
assign v$G2_13007_out0 = v$RD_6616_out0 && v$RM_12056_out0;
assign v$CARRY_5152_out0 = v$G2_12543_out0;
assign v$CARRY_5616_out0 = v$G2_13007_out0;
assign v$G1_7995_out0 = ((v$RD_6140_out0 && !v$RM_11580_out0) || (!v$RD_6140_out0) && v$RM_11580_out0);
assign v$G1_7997_out0 = ((v$RD_6142_out0 && !v$RM_11582_out0) || (!v$RD_6142_out0) && v$RM_11582_out0);
assign v$G1_8001_out0 = ((v$RD_6146_out0 && !v$RM_11586_out0) || (!v$RD_6146_out0) && v$RM_11586_out0);
assign v$G1_8003_out0 = ((v$RD_6148_out0 && !v$RM_11588_out0) || (!v$RD_6148_out0) && v$RM_11588_out0);
assign v$G1_8005_out0 = ((v$RD_6150_out0 && !v$RM_11590_out0) || (!v$RD_6150_out0) && v$RM_11590_out0);
assign v$G1_8008_out0 = ((v$RD_6153_out0 && !v$RM_11593_out0) || (!v$RD_6153_out0) && v$RM_11593_out0);
assign v$G1_8010_out0 = ((v$RD_6155_out0 && !v$RM_11595_out0) || (!v$RD_6155_out0) && v$RM_11595_out0);
assign v$G1_8012_out0 = ((v$RD_6157_out0 && !v$RM_11597_out0) || (!v$RD_6157_out0) && v$RM_11597_out0);
assign v$G1_8014_out0 = ((v$RD_6159_out0 && !v$RM_11599_out0) || (!v$RD_6159_out0) && v$RM_11599_out0);
assign v$G1_8016_out0 = ((v$RD_6161_out0 && !v$RM_11601_out0) || (!v$RD_6161_out0) && v$RM_11601_out0);
assign v$G1_8018_out0 = ((v$RD_6163_out0 && !v$RM_11603_out0) || (!v$RD_6163_out0) && v$RM_11603_out0);
assign v$G1_8020_out0 = ((v$RD_6165_out0 && !v$RM_11605_out0) || (!v$RD_6165_out0) && v$RM_11605_out0);
assign v$G1_8022_out0 = ((v$RD_6167_out0 && !v$RM_11607_out0) || (!v$RD_6167_out0) && v$RM_11607_out0);
assign v$G1_8024_out0 = ((v$RD_6169_out0 && !v$RM_11609_out0) || (!v$RD_6169_out0) && v$RM_11609_out0);
assign v$G1_8459_out0 = ((v$RD_6604_out0 && !v$RM_12044_out0) || (!v$RD_6604_out0) && v$RM_12044_out0);
assign v$G1_8461_out0 = ((v$RD_6606_out0 && !v$RM_12046_out0) || (!v$RD_6606_out0) && v$RM_12046_out0);
assign v$G1_8465_out0 = ((v$RD_6610_out0 && !v$RM_12050_out0) || (!v$RD_6610_out0) && v$RM_12050_out0);
assign v$G1_8467_out0 = ((v$RD_6612_out0 && !v$RM_12052_out0) || (!v$RD_6612_out0) && v$RM_12052_out0);
assign v$G1_8469_out0 = ((v$RD_6614_out0 && !v$RM_12054_out0) || (!v$RD_6614_out0) && v$RM_12054_out0);
assign v$G1_8472_out0 = ((v$RD_6617_out0 && !v$RM_12057_out0) || (!v$RD_6617_out0) && v$RM_12057_out0);
assign v$G1_8474_out0 = ((v$RD_6619_out0 && !v$RM_12059_out0) || (!v$RD_6619_out0) && v$RM_12059_out0);
assign v$G1_8476_out0 = ((v$RD_6621_out0 && !v$RM_12061_out0) || (!v$RD_6621_out0) && v$RM_12061_out0);
assign v$G1_8478_out0 = ((v$RD_6623_out0 && !v$RM_12063_out0) || (!v$RD_6623_out0) && v$RM_12063_out0);
assign v$G1_8480_out0 = ((v$RD_6625_out0 && !v$RM_12065_out0) || (!v$RD_6625_out0) && v$RM_12065_out0);
assign v$G1_8482_out0 = ((v$RD_6627_out0 && !v$RM_12067_out0) || (!v$RD_6627_out0) && v$RM_12067_out0);
assign v$G1_8484_out0 = ((v$RD_6629_out0 && !v$RM_12069_out0) || (!v$RD_6629_out0) && v$RM_12069_out0);
assign v$G1_8486_out0 = ((v$RD_6631_out0 && !v$RM_12071_out0) || (!v$RD_6631_out0) && v$RM_12071_out0);
assign v$G1_8488_out0 = ((v$RD_6633_out0 && !v$RM_12073_out0) || (!v$RD_6633_out0) && v$RM_12073_out0);
assign v$S_9153_out0 = v$G1_8007_out0;
assign v$S_9617_out0 = v$G1_8471_out0;
assign v$G2_12531_out0 = v$RD_6140_out0 && v$RM_11580_out0;
assign v$G2_12533_out0 = v$RD_6142_out0 && v$RM_11582_out0;
assign v$G2_12537_out0 = v$RD_6146_out0 && v$RM_11586_out0;
assign v$G2_12539_out0 = v$RD_6148_out0 && v$RM_11588_out0;
assign v$G2_12541_out0 = v$RD_6150_out0 && v$RM_11590_out0;
assign v$G2_12544_out0 = v$RD_6153_out0 && v$RM_11593_out0;
assign v$G2_12546_out0 = v$RD_6155_out0 && v$RM_11595_out0;
assign v$G2_12548_out0 = v$RD_6157_out0 && v$RM_11597_out0;
assign v$G2_12550_out0 = v$RD_6159_out0 && v$RM_11599_out0;
assign v$G2_12552_out0 = v$RD_6161_out0 && v$RM_11601_out0;
assign v$G2_12554_out0 = v$RD_6163_out0 && v$RM_11603_out0;
assign v$G2_12556_out0 = v$RD_6165_out0 && v$RM_11605_out0;
assign v$G2_12558_out0 = v$RD_6167_out0 && v$RM_11607_out0;
assign v$G2_12560_out0 = v$RD_6169_out0 && v$RM_11609_out0;
assign v$G2_12995_out0 = v$RD_6604_out0 && v$RM_12044_out0;
assign v$G2_12997_out0 = v$RD_6606_out0 && v$RM_12046_out0;
assign v$G2_13001_out0 = v$RD_6610_out0 && v$RM_12050_out0;
assign v$G2_13003_out0 = v$RD_6612_out0 && v$RM_12052_out0;
assign v$G2_13005_out0 = v$RD_6614_out0 && v$RM_12054_out0;
assign v$G2_13008_out0 = v$RD_6617_out0 && v$RM_12057_out0;
assign v$G2_13010_out0 = v$RD_6619_out0 && v$RM_12059_out0;
assign v$G2_13012_out0 = v$RD_6621_out0 && v$RM_12061_out0;
assign v$G2_13014_out0 = v$RD_6623_out0 && v$RM_12063_out0;
assign v$G2_13016_out0 = v$RD_6625_out0 && v$RM_12065_out0;
assign v$G2_13018_out0 = v$RD_6627_out0 && v$RM_12067_out0;
assign v$G2_13020_out0 = v$RD_6629_out0 && v$RM_12069_out0;
assign v$G2_13022_out0 = v$RD_6631_out0 && v$RM_12071_out0;
assign v$G2_13024_out0 = v$RD_6633_out0 && v$RM_12073_out0;
assign v$S_4674_out0 = v$S_9153_out0;
assign v$S_4689_out0 = v$S_9617_out0;
assign v$CARRY_5140_out0 = v$G2_12531_out0;
assign v$CARRY_5142_out0 = v$G2_12533_out0;
assign v$CARRY_5146_out0 = v$G2_12537_out0;
assign v$CARRY_5148_out0 = v$G2_12539_out0;
assign v$CARRY_5150_out0 = v$G2_12541_out0;
assign v$CARRY_5153_out0 = v$G2_12544_out0;
assign v$CARRY_5155_out0 = v$G2_12546_out0;
assign v$CARRY_5157_out0 = v$G2_12548_out0;
assign v$CARRY_5159_out0 = v$G2_12550_out0;
assign v$CARRY_5161_out0 = v$G2_12552_out0;
assign v$CARRY_5163_out0 = v$G2_12554_out0;
assign v$CARRY_5165_out0 = v$G2_12556_out0;
assign v$CARRY_5167_out0 = v$G2_12558_out0;
assign v$CARRY_5169_out0 = v$G2_12560_out0;
assign v$CARRY_5604_out0 = v$G2_12995_out0;
assign v$CARRY_5606_out0 = v$G2_12997_out0;
assign v$CARRY_5610_out0 = v$G2_13001_out0;
assign v$CARRY_5612_out0 = v$G2_13003_out0;
assign v$CARRY_5614_out0 = v$G2_13005_out0;
assign v$CARRY_5617_out0 = v$G2_13008_out0;
assign v$CARRY_5619_out0 = v$G2_13010_out0;
assign v$CARRY_5621_out0 = v$G2_13012_out0;
assign v$CARRY_5623_out0 = v$G2_13014_out0;
assign v$CARRY_5625_out0 = v$G2_13016_out0;
assign v$CARRY_5627_out0 = v$G2_13018_out0;
assign v$CARRY_5629_out0 = v$G2_13020_out0;
assign v$CARRY_5631_out0 = v$G2_13022_out0;
assign v$CARRY_5633_out0 = v$G2_13024_out0;
assign v$S_9141_out0 = v$G1_7995_out0;
assign v$S_9143_out0 = v$G1_7997_out0;
assign v$S_9147_out0 = v$G1_8001_out0;
assign v$S_9149_out0 = v$G1_8003_out0;
assign v$S_9151_out0 = v$G1_8005_out0;
assign v$S_9154_out0 = v$G1_8008_out0;
assign v$S_9156_out0 = v$G1_8010_out0;
assign v$S_9158_out0 = v$G1_8012_out0;
assign v$S_9160_out0 = v$G1_8014_out0;
assign v$S_9162_out0 = v$G1_8016_out0;
assign v$S_9164_out0 = v$G1_8018_out0;
assign v$S_9166_out0 = v$G1_8020_out0;
assign v$S_9168_out0 = v$G1_8022_out0;
assign v$S_9170_out0 = v$G1_8024_out0;
assign v$S_9605_out0 = v$G1_8459_out0;
assign v$S_9607_out0 = v$G1_8461_out0;
assign v$S_9611_out0 = v$G1_8465_out0;
assign v$S_9613_out0 = v$G1_8467_out0;
assign v$S_9615_out0 = v$G1_8469_out0;
assign v$S_9618_out0 = v$G1_8472_out0;
assign v$S_9620_out0 = v$G1_8474_out0;
assign v$S_9622_out0 = v$G1_8476_out0;
assign v$S_9624_out0 = v$G1_8478_out0;
assign v$S_9626_out0 = v$G1_8480_out0;
assign v$S_9628_out0 = v$G1_8482_out0;
assign v$S_9630_out0 = v$G1_8484_out0;
assign v$S_9632_out0 = v$G1_8486_out0;
assign v$S_9634_out0 = v$G1_8488_out0;
assign v$CIN_9950_out0 = v$CARRY_5152_out0;
assign v$CIN_10174_out0 = v$CARRY_5616_out0;
assign v$_43_out0 = { v$_636_out0,v$S_4674_out0 };
assign v$_44_out0 = { v$_637_out0,v$S_4689_out0 };
assign v$RD_6158_out0 = v$CIN_9950_out0;
assign v$RD_6622_out0 = v$CIN_10174_out0;
assign v$RM_11581_out0 = v$S_9141_out0;
assign v$RM_11583_out0 = v$S_9143_out0;
assign v$RM_11587_out0 = v$S_9147_out0;
assign v$RM_11589_out0 = v$S_9149_out0;
assign v$RM_11591_out0 = v$S_9151_out0;
assign v$RM_11594_out0 = v$S_9154_out0;
assign v$RM_11596_out0 = v$S_9156_out0;
assign v$RM_11598_out0 = v$S_9158_out0;
assign v$RM_11600_out0 = v$S_9160_out0;
assign v$RM_11602_out0 = v$S_9162_out0;
assign v$RM_11604_out0 = v$S_9164_out0;
assign v$RM_11606_out0 = v$S_9166_out0;
assign v$RM_11608_out0 = v$S_9168_out0;
assign v$RM_11610_out0 = v$S_9170_out0;
assign v$RM_12045_out0 = v$S_9605_out0;
assign v$RM_12047_out0 = v$S_9607_out0;
assign v$RM_12051_out0 = v$S_9611_out0;
assign v$RM_12053_out0 = v$S_9613_out0;
assign v$RM_12055_out0 = v$S_9615_out0;
assign v$RM_12058_out0 = v$S_9618_out0;
assign v$RM_12060_out0 = v$S_9620_out0;
assign v$RM_12062_out0 = v$S_9622_out0;
assign v$RM_12064_out0 = v$S_9624_out0;
assign v$RM_12066_out0 = v$S_9626_out0;
assign v$RM_12068_out0 = v$S_9628_out0;
assign v$RM_12070_out0 = v$S_9630_out0;
assign v$RM_12072_out0 = v$S_9632_out0;
assign v$RM_12074_out0 = v$S_9634_out0;
assign v$G1_8013_out0 = ((v$RD_6158_out0 && !v$RM_11598_out0) || (!v$RD_6158_out0) && v$RM_11598_out0);
assign v$G1_8477_out0 = ((v$RD_6622_out0 && !v$RM_12062_out0) || (!v$RD_6622_out0) && v$RM_12062_out0);
assign v$G2_12549_out0 = v$RD_6158_out0 && v$RM_11598_out0;
assign v$G2_13013_out0 = v$RD_6622_out0 && v$RM_12062_out0;
assign v$CARRY_5158_out0 = v$G2_12549_out0;
assign v$CARRY_5622_out0 = v$G2_13013_out0;
assign v$S_9159_out0 = v$G1_8013_out0;
assign v$S_9623_out0 = v$G1_8477_out0;
assign v$S_1361_out0 = v$S_9159_out0;
assign v$S_1585_out0 = v$S_9623_out0;
assign v$G1_4137_out0 = v$CARRY_5158_out0 || v$CARRY_5157_out0;
assign v$G1_4361_out0 = v$CARRY_5622_out0 || v$CARRY_5621_out0;
assign v$COUT_829_out0 = v$G1_4137_out0;
assign v$COUT_1053_out0 = v$G1_4361_out0;
assign v$CIN_9956_out0 = v$COUT_829_out0;
assign v$CIN_10180_out0 = v$COUT_1053_out0;
assign v$RD_6170_out0 = v$CIN_9956_out0;
assign v$RD_6634_out0 = v$CIN_10180_out0;
assign v$G1_8025_out0 = ((v$RD_6170_out0 && !v$RM_11610_out0) || (!v$RD_6170_out0) && v$RM_11610_out0);
assign v$G1_8489_out0 = ((v$RD_6634_out0 && !v$RM_12074_out0) || (!v$RD_6634_out0) && v$RM_12074_out0);
assign v$G2_12561_out0 = v$RD_6170_out0 && v$RM_11610_out0;
assign v$G2_13025_out0 = v$RD_6634_out0 && v$RM_12074_out0;
assign v$CARRY_5170_out0 = v$G2_12561_out0;
assign v$CARRY_5634_out0 = v$G2_13025_out0;
assign v$S_9171_out0 = v$G1_8025_out0;
assign v$S_9635_out0 = v$G1_8489_out0;
assign v$S_1367_out0 = v$S_9171_out0;
assign v$S_1591_out0 = v$S_9635_out0;
assign v$G1_4143_out0 = v$CARRY_5170_out0 || v$CARRY_5169_out0;
assign v$G1_4367_out0 = v$CARRY_5634_out0 || v$CARRY_5633_out0;
assign v$COUT_835_out0 = v$G1_4143_out0;
assign v$COUT_1059_out0 = v$G1_4367_out0;
assign v$_4791_out0 = { v$S_1361_out0,v$S_1367_out0 };
assign v$_4806_out0 = { v$S_1585_out0,v$S_1591_out0 };
assign v$CIN_9951_out0 = v$COUT_835_out0;
assign v$CIN_10175_out0 = v$COUT_1059_out0;
assign v$RD_6160_out0 = v$CIN_9951_out0;
assign v$RD_6624_out0 = v$CIN_10175_out0;
assign v$G1_8015_out0 = ((v$RD_6160_out0 && !v$RM_11600_out0) || (!v$RD_6160_out0) && v$RM_11600_out0);
assign v$G1_8479_out0 = ((v$RD_6624_out0 && !v$RM_12064_out0) || (!v$RD_6624_out0) && v$RM_12064_out0);
assign v$G2_12551_out0 = v$RD_6160_out0 && v$RM_11600_out0;
assign v$G2_13015_out0 = v$RD_6624_out0 && v$RM_12064_out0;
assign v$CARRY_5160_out0 = v$G2_12551_out0;
assign v$CARRY_5624_out0 = v$G2_13015_out0;
assign v$S_9161_out0 = v$G1_8015_out0;
assign v$S_9625_out0 = v$G1_8479_out0;
assign v$S_1362_out0 = v$S_9161_out0;
assign v$S_1586_out0 = v$S_9625_out0;
assign v$G1_4138_out0 = v$CARRY_5160_out0 || v$CARRY_5159_out0;
assign v$G1_4362_out0 = v$CARRY_5624_out0 || v$CARRY_5623_out0;
assign v$COUT_830_out0 = v$G1_4138_out0;
assign v$COUT_1054_out0 = v$G1_4362_out0;
assign v$_2561_out0 = { v$_4791_out0,v$S_1362_out0 };
assign v$_2576_out0 = { v$_4806_out0,v$S_1586_out0 };
assign v$CIN_9946_out0 = v$COUT_830_out0;
assign v$CIN_10170_out0 = v$COUT_1054_out0;
assign v$RD_6149_out0 = v$CIN_9946_out0;
assign v$RD_6613_out0 = v$CIN_10170_out0;
assign v$G1_8004_out0 = ((v$RD_6149_out0 && !v$RM_11589_out0) || (!v$RD_6149_out0) && v$RM_11589_out0);
assign v$G1_8468_out0 = ((v$RD_6613_out0 && !v$RM_12053_out0) || (!v$RD_6613_out0) && v$RM_12053_out0);
assign v$G2_12540_out0 = v$RD_6149_out0 && v$RM_11589_out0;
assign v$G2_13004_out0 = v$RD_6613_out0 && v$RM_12053_out0;
assign v$CARRY_5149_out0 = v$G2_12540_out0;
assign v$CARRY_5613_out0 = v$G2_13004_out0;
assign v$S_9150_out0 = v$G1_8004_out0;
assign v$S_9614_out0 = v$G1_8468_out0;
assign v$S_1357_out0 = v$S_9150_out0;
assign v$S_1581_out0 = v$S_9614_out0;
assign v$G1_4133_out0 = v$CARRY_5149_out0 || v$CARRY_5148_out0;
assign v$G1_4357_out0 = v$CARRY_5613_out0 || v$CARRY_5612_out0;
assign v$COUT_825_out0 = v$G1_4133_out0;
assign v$COUT_1049_out0 = v$G1_4357_out0;
assign v$_7041_out0 = { v$_2561_out0,v$S_1357_out0 };
assign v$_7056_out0 = { v$_2576_out0,v$S_1581_out0 };
assign v$CIN_9945_out0 = v$COUT_825_out0;
assign v$CIN_10169_out0 = v$COUT_1049_out0;
assign v$RD_6147_out0 = v$CIN_9945_out0;
assign v$RD_6611_out0 = v$CIN_10169_out0;
assign v$G1_8002_out0 = ((v$RD_6147_out0 && !v$RM_11587_out0) || (!v$RD_6147_out0) && v$RM_11587_out0);
assign v$G1_8466_out0 = ((v$RD_6611_out0 && !v$RM_12051_out0) || (!v$RD_6611_out0) && v$RM_12051_out0);
assign v$G2_12538_out0 = v$RD_6147_out0 && v$RM_11587_out0;
assign v$G2_13002_out0 = v$RD_6611_out0 && v$RM_12051_out0;
assign v$CARRY_5147_out0 = v$G2_12538_out0;
assign v$CARRY_5611_out0 = v$G2_13002_out0;
assign v$S_9148_out0 = v$G1_8002_out0;
assign v$S_9612_out0 = v$G1_8466_out0;
assign v$S_1356_out0 = v$S_9148_out0;
assign v$S_1580_out0 = v$S_9612_out0;
assign v$G1_4132_out0 = v$CARRY_5147_out0 || v$CARRY_5146_out0;
assign v$G1_4356_out0 = v$CARRY_5611_out0 || v$CARRY_5610_out0;
assign v$COUT_824_out0 = v$G1_4132_out0;
assign v$COUT_1048_out0 = v$G1_4356_out0;
assign v$_13527_out0 = { v$_7041_out0,v$S_1356_out0 };
assign v$_13542_out0 = { v$_7056_out0,v$S_1580_out0 };
assign v$CIN_9952_out0 = v$COUT_824_out0;
assign v$CIN_10176_out0 = v$COUT_1048_out0;
assign v$RD_6162_out0 = v$CIN_9952_out0;
assign v$RD_6626_out0 = v$CIN_10176_out0;
assign v$G1_8017_out0 = ((v$RD_6162_out0 && !v$RM_11602_out0) || (!v$RD_6162_out0) && v$RM_11602_out0);
assign v$G1_8481_out0 = ((v$RD_6626_out0 && !v$RM_12066_out0) || (!v$RD_6626_out0) && v$RM_12066_out0);
assign v$G2_12553_out0 = v$RD_6162_out0 && v$RM_11602_out0;
assign v$G2_13017_out0 = v$RD_6626_out0 && v$RM_12066_out0;
assign v$CARRY_5162_out0 = v$G2_12553_out0;
assign v$CARRY_5626_out0 = v$G2_13017_out0;
assign v$S_9163_out0 = v$G1_8017_out0;
assign v$S_9627_out0 = v$G1_8481_out0;
assign v$S_1363_out0 = v$S_9163_out0;
assign v$S_1587_out0 = v$S_9627_out0;
assign v$G1_4139_out0 = v$CARRY_5162_out0 || v$CARRY_5161_out0;
assign v$G1_4363_out0 = v$CARRY_5626_out0 || v$CARRY_5625_out0;
assign v$COUT_831_out0 = v$G1_4139_out0;
assign v$COUT_1055_out0 = v$G1_4363_out0;
assign v$_3320_out0 = { v$_13527_out0,v$S_1363_out0 };
assign v$_3335_out0 = { v$_13542_out0,v$S_1587_out0 };
assign v$CIN_9953_out0 = v$COUT_831_out0;
assign v$CIN_10177_out0 = v$COUT_1055_out0;
assign v$RD_6164_out0 = v$CIN_9953_out0;
assign v$RD_6628_out0 = v$CIN_10177_out0;
assign v$G1_8019_out0 = ((v$RD_6164_out0 && !v$RM_11604_out0) || (!v$RD_6164_out0) && v$RM_11604_out0);
assign v$G1_8483_out0 = ((v$RD_6628_out0 && !v$RM_12068_out0) || (!v$RD_6628_out0) && v$RM_12068_out0);
assign v$G2_12555_out0 = v$RD_6164_out0 && v$RM_11604_out0;
assign v$G2_13019_out0 = v$RD_6628_out0 && v$RM_12068_out0;
assign v$CARRY_5164_out0 = v$G2_12555_out0;
assign v$CARRY_5628_out0 = v$G2_13019_out0;
assign v$S_9165_out0 = v$G1_8019_out0;
assign v$S_9629_out0 = v$G1_8483_out0;
assign v$S_1364_out0 = v$S_9165_out0;
assign v$S_1588_out0 = v$S_9629_out0;
assign v$G1_4140_out0 = v$CARRY_5164_out0 || v$CARRY_5163_out0;
assign v$G1_4364_out0 = v$CARRY_5628_out0 || v$CARRY_5627_out0;
assign v$COUT_832_out0 = v$G1_4140_out0;
assign v$COUT_1056_out0 = v$G1_4364_out0;
assign v$_7156_out0 = { v$_3320_out0,v$S_1364_out0 };
assign v$_7171_out0 = { v$_3335_out0,v$S_1588_out0 };
assign v$CIN_9955_out0 = v$COUT_832_out0;
assign v$CIN_10179_out0 = v$COUT_1056_out0;
assign v$RD_6168_out0 = v$CIN_9955_out0;
assign v$RD_6632_out0 = v$CIN_10179_out0;
assign v$G1_8023_out0 = ((v$RD_6168_out0 && !v$RM_11608_out0) || (!v$RD_6168_out0) && v$RM_11608_out0);
assign v$G1_8487_out0 = ((v$RD_6632_out0 && !v$RM_12072_out0) || (!v$RD_6632_out0) && v$RM_12072_out0);
assign v$G2_12559_out0 = v$RD_6168_out0 && v$RM_11608_out0;
assign v$G2_13023_out0 = v$RD_6632_out0 && v$RM_12072_out0;
assign v$CARRY_5168_out0 = v$G2_12559_out0;
assign v$CARRY_5632_out0 = v$G2_13023_out0;
assign v$S_9169_out0 = v$G1_8023_out0;
assign v$S_9633_out0 = v$G1_8487_out0;
assign v$S_1366_out0 = v$S_9169_out0;
assign v$S_1590_out0 = v$S_9633_out0;
assign v$G1_4142_out0 = v$CARRY_5168_out0 || v$CARRY_5167_out0;
assign v$G1_4366_out0 = v$CARRY_5632_out0 || v$CARRY_5631_out0;
assign v$COUT_834_out0 = v$G1_4142_out0;
assign v$COUT_1058_out0 = v$G1_4366_out0;
assign v$_4758_out0 = { v$_7156_out0,v$S_1366_out0 };
assign v$_4773_out0 = { v$_7171_out0,v$S_1590_out0 };
assign v$CIN_9948_out0 = v$COUT_834_out0;
assign v$CIN_10172_out0 = v$COUT_1058_out0;
assign v$RD_6154_out0 = v$CIN_9948_out0;
assign v$RD_6618_out0 = v$CIN_10172_out0;
assign v$G1_8009_out0 = ((v$RD_6154_out0 && !v$RM_11594_out0) || (!v$RD_6154_out0) && v$RM_11594_out0);
assign v$G1_8473_out0 = ((v$RD_6618_out0 && !v$RM_12058_out0) || (!v$RD_6618_out0) && v$RM_12058_out0);
assign v$G2_12545_out0 = v$RD_6154_out0 && v$RM_11594_out0;
assign v$G2_13009_out0 = v$RD_6618_out0 && v$RM_12058_out0;
assign v$CARRY_5154_out0 = v$G2_12545_out0;
assign v$CARRY_5618_out0 = v$G2_13009_out0;
assign v$S_9155_out0 = v$G1_8009_out0;
assign v$S_9619_out0 = v$G1_8473_out0;
assign v$S_1359_out0 = v$S_9155_out0;
assign v$S_1583_out0 = v$S_9619_out0;
assign v$G1_4135_out0 = v$CARRY_5154_out0 || v$CARRY_5153_out0;
assign v$G1_4359_out0 = v$CARRY_5618_out0 || v$CARRY_5617_out0;
assign v$COUT_827_out0 = v$G1_4135_out0;
assign v$COUT_1051_out0 = v$G1_4359_out0;
assign v$_6935_out0 = { v$_4758_out0,v$S_1359_out0 };
assign v$_6950_out0 = { v$_4773_out0,v$S_1583_out0 };
assign v$CIN_9949_out0 = v$COUT_827_out0;
assign v$CIN_10173_out0 = v$COUT_1051_out0;
assign v$RD_6156_out0 = v$CIN_9949_out0;
assign v$RD_6620_out0 = v$CIN_10173_out0;
assign v$G1_8011_out0 = ((v$RD_6156_out0 && !v$RM_11596_out0) || (!v$RD_6156_out0) && v$RM_11596_out0);
assign v$G1_8475_out0 = ((v$RD_6620_out0 && !v$RM_12060_out0) || (!v$RD_6620_out0) && v$RM_12060_out0);
assign v$G2_12547_out0 = v$RD_6156_out0 && v$RM_11596_out0;
assign v$G2_13011_out0 = v$RD_6620_out0 && v$RM_12060_out0;
assign v$CARRY_5156_out0 = v$G2_12547_out0;
assign v$CARRY_5620_out0 = v$G2_13011_out0;
assign v$S_9157_out0 = v$G1_8011_out0;
assign v$S_9621_out0 = v$G1_8475_out0;
assign v$S_1360_out0 = v$S_9157_out0;
assign v$S_1584_out0 = v$S_9621_out0;
assign v$G1_4136_out0 = v$CARRY_5156_out0 || v$CARRY_5155_out0;
assign v$G1_4360_out0 = v$CARRY_5620_out0 || v$CARRY_5619_out0;
assign v$COUT_828_out0 = v$G1_4136_out0;
assign v$COUT_1052_out0 = v$G1_4360_out0;
assign v$_5811_out0 = { v$_6935_out0,v$S_1360_out0 };
assign v$_5826_out0 = { v$_6950_out0,v$S_1584_out0 };
assign v$CIN_9954_out0 = v$COUT_828_out0;
assign v$CIN_10178_out0 = v$COUT_1052_out0;
assign v$RD_6166_out0 = v$CIN_9954_out0;
assign v$RD_6630_out0 = v$CIN_10178_out0;
assign v$G1_8021_out0 = ((v$RD_6166_out0 && !v$RM_11606_out0) || (!v$RD_6166_out0) && v$RM_11606_out0);
assign v$G1_8485_out0 = ((v$RD_6630_out0 && !v$RM_12070_out0) || (!v$RD_6630_out0) && v$RM_12070_out0);
assign v$G2_12557_out0 = v$RD_6166_out0 && v$RM_11606_out0;
assign v$G2_13021_out0 = v$RD_6630_out0 && v$RM_12070_out0;
assign v$CARRY_5166_out0 = v$G2_12557_out0;
assign v$CARRY_5630_out0 = v$G2_13021_out0;
assign v$S_9167_out0 = v$G1_8021_out0;
assign v$S_9631_out0 = v$G1_8485_out0;
assign v$S_1365_out0 = v$S_9167_out0;
assign v$S_1589_out0 = v$S_9631_out0;
assign v$G1_4141_out0 = v$CARRY_5166_out0 || v$CARRY_5165_out0;
assign v$G1_4365_out0 = v$CARRY_5630_out0 || v$CARRY_5629_out0;
assign v$COUT_833_out0 = v$G1_4141_out0;
assign v$COUT_1057_out0 = v$G1_4365_out0;
assign v$_2035_out0 = { v$_5811_out0,v$S_1365_out0 };
assign v$_2050_out0 = { v$_5826_out0,v$S_1589_out0 };
assign v$CIN_9942_out0 = v$COUT_833_out0;
assign v$CIN_10166_out0 = v$COUT_1057_out0;
assign v$RD_6141_out0 = v$CIN_9942_out0;
assign v$RD_6605_out0 = v$CIN_10166_out0;
assign v$G1_7996_out0 = ((v$RD_6141_out0 && !v$RM_11581_out0) || (!v$RD_6141_out0) && v$RM_11581_out0);
assign v$G1_8460_out0 = ((v$RD_6605_out0 && !v$RM_12045_out0) || (!v$RD_6605_out0) && v$RM_12045_out0);
assign v$G2_12532_out0 = v$RD_6141_out0 && v$RM_11581_out0;
assign v$G2_12996_out0 = v$RD_6605_out0 && v$RM_12045_out0;
assign v$CARRY_5141_out0 = v$G2_12532_out0;
assign v$CARRY_5605_out0 = v$G2_12996_out0;
assign v$S_9142_out0 = v$G1_7996_out0;
assign v$S_9606_out0 = v$G1_8460_out0;
assign v$S_1353_out0 = v$S_9142_out0;
assign v$S_1577_out0 = v$S_9606_out0;
assign v$G1_4129_out0 = v$CARRY_5141_out0 || v$CARRY_5140_out0;
assign v$G1_4353_out0 = v$CARRY_5605_out0 || v$CARRY_5604_out0;
assign v$COUT_821_out0 = v$G1_4129_out0;
assign v$COUT_1045_out0 = v$G1_4353_out0;
assign v$_2802_out0 = { v$_2035_out0,v$S_1353_out0 };
assign v$_2817_out0 = { v$_2050_out0,v$S_1577_out0 };
assign v$CIN_9947_out0 = v$COUT_821_out0;
assign v$CIN_10171_out0 = v$COUT_1045_out0;
assign v$RD_6151_out0 = v$CIN_9947_out0;
assign v$RD_6615_out0 = v$CIN_10171_out0;
assign v$G1_8006_out0 = ((v$RD_6151_out0 && !v$RM_11591_out0) || (!v$RD_6151_out0) && v$RM_11591_out0);
assign v$G1_8470_out0 = ((v$RD_6615_out0 && !v$RM_12055_out0) || (!v$RD_6615_out0) && v$RM_12055_out0);
assign v$G2_12542_out0 = v$RD_6151_out0 && v$RM_11591_out0;
assign v$G2_13006_out0 = v$RD_6615_out0 && v$RM_12055_out0;
assign v$CARRY_5151_out0 = v$G2_12542_out0;
assign v$CARRY_5615_out0 = v$G2_13006_out0;
assign v$S_9152_out0 = v$G1_8006_out0;
assign v$S_9616_out0 = v$G1_8470_out0;
assign v$S_1358_out0 = v$S_9152_out0;
assign v$S_1582_out0 = v$S_9616_out0;
assign v$G1_4134_out0 = v$CARRY_5151_out0 || v$CARRY_5150_out0;
assign v$G1_4358_out0 = v$CARRY_5615_out0 || v$CARRY_5614_out0;
assign v$COUT_826_out0 = v$G1_4134_out0;
assign v$COUT_1050_out0 = v$G1_4358_out0;
assign v$_1834_out0 = { v$_2802_out0,v$S_1358_out0 };
assign v$_1849_out0 = { v$_2817_out0,v$S_1582_out0 };
assign v$CIN_9943_out0 = v$COUT_826_out0;
assign v$CIN_10167_out0 = v$COUT_1050_out0;
assign v$RD_6143_out0 = v$CIN_9943_out0;
assign v$RD_6607_out0 = v$CIN_10167_out0;
assign v$G1_7998_out0 = ((v$RD_6143_out0 && !v$RM_11583_out0) || (!v$RD_6143_out0) && v$RM_11583_out0);
assign v$G1_8462_out0 = ((v$RD_6607_out0 && !v$RM_12047_out0) || (!v$RD_6607_out0) && v$RM_12047_out0);
assign v$G2_12534_out0 = v$RD_6143_out0 && v$RM_11583_out0;
assign v$G2_12998_out0 = v$RD_6607_out0 && v$RM_12047_out0;
assign v$CARRY_5143_out0 = v$G2_12534_out0;
assign v$CARRY_5607_out0 = v$G2_12998_out0;
assign v$S_9144_out0 = v$G1_7998_out0;
assign v$S_9608_out0 = v$G1_8462_out0;
assign v$S_1354_out0 = v$S_9144_out0;
assign v$S_1578_out0 = v$S_9608_out0;
assign v$G1_4130_out0 = v$CARRY_5143_out0 || v$CARRY_5142_out0;
assign v$G1_4354_out0 = v$CARRY_5607_out0 || v$CARRY_5606_out0;
assign v$COUT_822_out0 = v$G1_4130_out0;
assign v$COUT_1046_out0 = v$G1_4354_out0;
assign v$_4558_out0 = { v$_1834_out0,v$S_1354_out0 };
assign v$_4573_out0 = { v$_1849_out0,v$S_1578_out0 };
assign v$RM_3491_out0 = v$COUT_822_out0;
assign v$RM_3715_out0 = v$COUT_1046_out0;
assign v$RM_11584_out0 = v$RM_3491_out0;
assign v$RM_12048_out0 = v$RM_3715_out0;
assign v$G1_7999_out0 = ((v$RD_6144_out0 && !v$RM_11584_out0) || (!v$RD_6144_out0) && v$RM_11584_out0);
assign v$G1_8463_out0 = ((v$RD_6608_out0 && !v$RM_12048_out0) || (!v$RD_6608_out0) && v$RM_12048_out0);
assign v$G2_12535_out0 = v$RD_6144_out0 && v$RM_11584_out0;
assign v$G2_12999_out0 = v$RD_6608_out0 && v$RM_12048_out0;
assign v$CARRY_5144_out0 = v$G2_12535_out0;
assign v$CARRY_5608_out0 = v$G2_12999_out0;
assign v$S_9145_out0 = v$G1_7999_out0;
assign v$S_9609_out0 = v$G1_8463_out0;
assign v$RM_11585_out0 = v$S_9145_out0;
assign v$RM_12049_out0 = v$S_9609_out0;
assign v$G1_8000_out0 = ((v$RD_6145_out0 && !v$RM_11585_out0) || (!v$RD_6145_out0) && v$RM_11585_out0);
assign v$G1_8464_out0 = ((v$RD_6609_out0 && !v$RM_12049_out0) || (!v$RD_6609_out0) && v$RM_12049_out0);
assign v$G2_12536_out0 = v$RD_6145_out0 && v$RM_11585_out0;
assign v$G2_13000_out0 = v$RD_6609_out0 && v$RM_12049_out0;
assign v$CARRY_5145_out0 = v$G2_12536_out0;
assign v$CARRY_5609_out0 = v$G2_13000_out0;
assign v$S_9146_out0 = v$G1_8000_out0;
assign v$S_9610_out0 = v$G1_8464_out0;
assign v$S_1355_out0 = v$S_9146_out0;
assign v$S_1579_out0 = v$S_9610_out0;
assign v$G1_4131_out0 = v$CARRY_5145_out0 || v$CARRY_5144_out0;
assign v$G1_4355_out0 = v$CARRY_5609_out0 || v$CARRY_5608_out0;
assign v$COUT_823_out0 = v$G1_4131_out0;
assign v$COUT_1047_out0 = v$G1_4355_out0;
assign v$_10660_out0 = { v$_4558_out0,v$S_1355_out0 };
assign v$_10675_out0 = { v$_4573_out0,v$S_1579_out0 };
assign v$_10955_out0 = { v$_10660_out0,v$COUT_823_out0 };
assign v$_10970_out0 = { v$_10675_out0,v$COUT_1047_out0 };
assign v$COUT_10925_out0 = v$_10955_out0;
assign v$COUT_10940_out0 = v$_10970_out0;
assign v$CIN_2369_out0 = v$COUT_10925_out0;
assign v$CIN_2384_out0 = v$COUT_10940_out0;
assign v$_482_out0 = v$CIN_2369_out0[8:8];
assign v$_497_out0 = v$CIN_2384_out0[8:8];
assign v$_1787_out0 = v$CIN_2369_out0[6:6];
assign v$_1802_out0 = v$CIN_2384_out0[6:6];
assign v$_2169_out0 = v$CIN_2369_out0[3:3];
assign v$_2184_out0 = v$CIN_2384_out0[3:3];
assign v$_2208_out0 = v$CIN_2369_out0[15:15];
assign v$_2222_out0 = v$CIN_2384_out0[15:15];
assign v$_2516_out0 = v$CIN_2369_out0[0:0];
assign v$_2531_out0 = v$CIN_2384_out0[0:0];
assign v$_3065_out0 = v$CIN_2369_out0[9:9];
assign v$_3080_out0 = v$CIN_2384_out0[9:9];
assign v$_3099_out0 = v$CIN_2369_out0[2:2];
assign v$_3114_out0 = v$CIN_2384_out0[2:2];
assign v$_3153_out0 = v$CIN_2369_out0[7:7];
assign v$_3168_out0 = v$CIN_2384_out0[7:7];
assign v$_3837_out0 = v$CIN_2369_out0[1:1];
assign v$_3852_out0 = v$CIN_2384_out0[1:1];
assign v$_3875_out0 = v$CIN_2369_out0[10:10];
assign v$_3890_out0 = v$CIN_2384_out0[10:10];
assign v$_6814_out0 = v$CIN_2369_out0[11:11];
assign v$_6829_out0 = v$CIN_2384_out0[11:11];
assign v$_7658_out0 = v$CIN_2369_out0[12:12];
assign v$_7673_out0 = v$CIN_2384_out0[12:12];
assign v$_8713_out0 = v$CIN_2369_out0[13:13];
assign v$_8728_out0 = v$CIN_2384_out0[13:13];
assign v$_8783_out0 = v$CIN_2369_out0[14:14];
assign v$_8798_out0 = v$CIN_2384_out0[14:14];
assign v$_10733_out0 = v$CIN_2369_out0[5:5];
assign v$_10748_out0 = v$CIN_2384_out0[5:5];
assign v$_13462_out0 = v$CIN_2369_out0[4:4];
assign v$_13477_out0 = v$CIN_2384_out0[4:4];
assign v$RM_3564_out0 = v$_7658_out0;
assign v$RM_3565_out0 = v$_8783_out0;
assign v$RM_3567_out0 = v$_10733_out0;
assign v$RM_3568_out0 = v$_13462_out0;
assign v$RM_3569_out0 = v$_8713_out0;
assign v$RM_3570_out0 = v$_3065_out0;
assign v$RM_3571_out0 = v$_3875_out0;
assign v$RM_3572_out0 = v$_3837_out0;
assign v$RM_3573_out0 = v$_2169_out0;
assign v$RM_3574_out0 = v$_1787_out0;
assign v$RM_3575_out0 = v$_3153_out0;
assign v$RM_3576_out0 = v$_6814_out0;
assign v$RM_3577_out0 = v$_482_out0;
assign v$RM_3578_out0 = v$_3099_out0;
assign v$RM_3788_out0 = v$_7673_out0;
assign v$RM_3789_out0 = v$_8798_out0;
assign v$RM_3791_out0 = v$_10748_out0;
assign v$RM_3792_out0 = v$_13477_out0;
assign v$RM_3793_out0 = v$_8728_out0;
assign v$RM_3794_out0 = v$_3080_out0;
assign v$RM_3795_out0 = v$_3890_out0;
assign v$RM_3796_out0 = v$_3852_out0;
assign v$RM_3797_out0 = v$_2184_out0;
assign v$RM_3798_out0 = v$_1802_out0;
assign v$RM_3799_out0 = v$_3168_out0;
assign v$RM_3800_out0 = v$_6829_out0;
assign v$RM_3801_out0 = v$_497_out0;
assign v$RM_3802_out0 = v$_3114_out0;
assign v$CIN_10019_out0 = v$_2208_out0;
assign v$CIN_10243_out0 = v$_2222_out0;
assign v$RM_11747_out0 = v$_2516_out0;
assign v$RM_12211_out0 = v$_2531_out0;
assign v$RD_6300_out0 = v$CIN_10019_out0;
assign v$RD_6764_out0 = v$CIN_10243_out0;
assign v$G1_8162_out0 = ((v$RD_6307_out0 && !v$RM_11747_out0) || (!v$RD_6307_out0) && v$RM_11747_out0);
assign v$G1_8626_out0 = ((v$RD_6771_out0 && !v$RM_12211_out0) || (!v$RD_6771_out0) && v$RM_12211_out0);
assign v$RM_11735_out0 = v$RM_3564_out0;
assign v$RM_11737_out0 = v$RM_3565_out0;
assign v$RM_11741_out0 = v$RM_3567_out0;
assign v$RM_11743_out0 = v$RM_3568_out0;
assign v$RM_11745_out0 = v$RM_3569_out0;
assign v$RM_11748_out0 = v$RM_3570_out0;
assign v$RM_11750_out0 = v$RM_3571_out0;
assign v$RM_11752_out0 = v$RM_3572_out0;
assign v$RM_11754_out0 = v$RM_3573_out0;
assign v$RM_11756_out0 = v$RM_3574_out0;
assign v$RM_11758_out0 = v$RM_3575_out0;
assign v$RM_11760_out0 = v$RM_3576_out0;
assign v$RM_11762_out0 = v$RM_3577_out0;
assign v$RM_11764_out0 = v$RM_3578_out0;
assign v$RM_12199_out0 = v$RM_3788_out0;
assign v$RM_12201_out0 = v$RM_3789_out0;
assign v$RM_12205_out0 = v$RM_3791_out0;
assign v$RM_12207_out0 = v$RM_3792_out0;
assign v$RM_12209_out0 = v$RM_3793_out0;
assign v$RM_12212_out0 = v$RM_3794_out0;
assign v$RM_12214_out0 = v$RM_3795_out0;
assign v$RM_12216_out0 = v$RM_3796_out0;
assign v$RM_12218_out0 = v$RM_3797_out0;
assign v$RM_12220_out0 = v$RM_3798_out0;
assign v$RM_12222_out0 = v$RM_3799_out0;
assign v$RM_12224_out0 = v$RM_3800_out0;
assign v$RM_12226_out0 = v$RM_3801_out0;
assign v$RM_12228_out0 = v$RM_3802_out0;
assign v$G2_12698_out0 = v$RD_6307_out0 && v$RM_11747_out0;
assign v$G2_13162_out0 = v$RD_6771_out0 && v$RM_12211_out0;
assign v$CARRY_5307_out0 = v$G2_12698_out0;
assign v$CARRY_5771_out0 = v$G2_13162_out0;
assign v$G1_8150_out0 = ((v$RD_6295_out0 && !v$RM_11735_out0) || (!v$RD_6295_out0) && v$RM_11735_out0);
assign v$G1_8152_out0 = ((v$RD_6297_out0 && !v$RM_11737_out0) || (!v$RD_6297_out0) && v$RM_11737_out0);
assign v$G1_8156_out0 = ((v$RD_6301_out0 && !v$RM_11741_out0) || (!v$RD_6301_out0) && v$RM_11741_out0);
assign v$G1_8158_out0 = ((v$RD_6303_out0 && !v$RM_11743_out0) || (!v$RD_6303_out0) && v$RM_11743_out0);
assign v$G1_8160_out0 = ((v$RD_6305_out0 && !v$RM_11745_out0) || (!v$RD_6305_out0) && v$RM_11745_out0);
assign v$G1_8163_out0 = ((v$RD_6308_out0 && !v$RM_11748_out0) || (!v$RD_6308_out0) && v$RM_11748_out0);
assign v$G1_8165_out0 = ((v$RD_6310_out0 && !v$RM_11750_out0) || (!v$RD_6310_out0) && v$RM_11750_out0);
assign v$G1_8167_out0 = ((v$RD_6312_out0 && !v$RM_11752_out0) || (!v$RD_6312_out0) && v$RM_11752_out0);
assign v$G1_8169_out0 = ((v$RD_6314_out0 && !v$RM_11754_out0) || (!v$RD_6314_out0) && v$RM_11754_out0);
assign v$G1_8171_out0 = ((v$RD_6316_out0 && !v$RM_11756_out0) || (!v$RD_6316_out0) && v$RM_11756_out0);
assign v$G1_8173_out0 = ((v$RD_6318_out0 && !v$RM_11758_out0) || (!v$RD_6318_out0) && v$RM_11758_out0);
assign v$G1_8175_out0 = ((v$RD_6320_out0 && !v$RM_11760_out0) || (!v$RD_6320_out0) && v$RM_11760_out0);
assign v$G1_8177_out0 = ((v$RD_6322_out0 && !v$RM_11762_out0) || (!v$RD_6322_out0) && v$RM_11762_out0);
assign v$G1_8179_out0 = ((v$RD_6324_out0 && !v$RM_11764_out0) || (!v$RD_6324_out0) && v$RM_11764_out0);
assign v$G1_8614_out0 = ((v$RD_6759_out0 && !v$RM_12199_out0) || (!v$RD_6759_out0) && v$RM_12199_out0);
assign v$G1_8616_out0 = ((v$RD_6761_out0 && !v$RM_12201_out0) || (!v$RD_6761_out0) && v$RM_12201_out0);
assign v$G1_8620_out0 = ((v$RD_6765_out0 && !v$RM_12205_out0) || (!v$RD_6765_out0) && v$RM_12205_out0);
assign v$G1_8622_out0 = ((v$RD_6767_out0 && !v$RM_12207_out0) || (!v$RD_6767_out0) && v$RM_12207_out0);
assign v$G1_8624_out0 = ((v$RD_6769_out0 && !v$RM_12209_out0) || (!v$RD_6769_out0) && v$RM_12209_out0);
assign v$G1_8627_out0 = ((v$RD_6772_out0 && !v$RM_12212_out0) || (!v$RD_6772_out0) && v$RM_12212_out0);
assign v$G1_8629_out0 = ((v$RD_6774_out0 && !v$RM_12214_out0) || (!v$RD_6774_out0) && v$RM_12214_out0);
assign v$G1_8631_out0 = ((v$RD_6776_out0 && !v$RM_12216_out0) || (!v$RD_6776_out0) && v$RM_12216_out0);
assign v$G1_8633_out0 = ((v$RD_6778_out0 && !v$RM_12218_out0) || (!v$RD_6778_out0) && v$RM_12218_out0);
assign v$G1_8635_out0 = ((v$RD_6780_out0 && !v$RM_12220_out0) || (!v$RD_6780_out0) && v$RM_12220_out0);
assign v$G1_8637_out0 = ((v$RD_6782_out0 && !v$RM_12222_out0) || (!v$RD_6782_out0) && v$RM_12222_out0);
assign v$G1_8639_out0 = ((v$RD_6784_out0 && !v$RM_12224_out0) || (!v$RD_6784_out0) && v$RM_12224_out0);
assign v$G1_8641_out0 = ((v$RD_6786_out0 && !v$RM_12226_out0) || (!v$RD_6786_out0) && v$RM_12226_out0);
assign v$G1_8643_out0 = ((v$RD_6788_out0 && !v$RM_12228_out0) || (!v$RD_6788_out0) && v$RM_12228_out0);
assign v$S_9308_out0 = v$G1_8162_out0;
assign v$S_9772_out0 = v$G1_8626_out0;
assign v$G2_12686_out0 = v$RD_6295_out0 && v$RM_11735_out0;
assign v$G2_12688_out0 = v$RD_6297_out0 && v$RM_11737_out0;
assign v$G2_12692_out0 = v$RD_6301_out0 && v$RM_11741_out0;
assign v$G2_12694_out0 = v$RD_6303_out0 && v$RM_11743_out0;
assign v$G2_12696_out0 = v$RD_6305_out0 && v$RM_11745_out0;
assign v$G2_12699_out0 = v$RD_6308_out0 && v$RM_11748_out0;
assign v$G2_12701_out0 = v$RD_6310_out0 && v$RM_11750_out0;
assign v$G2_12703_out0 = v$RD_6312_out0 && v$RM_11752_out0;
assign v$G2_12705_out0 = v$RD_6314_out0 && v$RM_11754_out0;
assign v$G2_12707_out0 = v$RD_6316_out0 && v$RM_11756_out0;
assign v$G2_12709_out0 = v$RD_6318_out0 && v$RM_11758_out0;
assign v$G2_12711_out0 = v$RD_6320_out0 && v$RM_11760_out0;
assign v$G2_12713_out0 = v$RD_6322_out0 && v$RM_11762_out0;
assign v$G2_12715_out0 = v$RD_6324_out0 && v$RM_11764_out0;
assign v$G2_13150_out0 = v$RD_6759_out0 && v$RM_12199_out0;
assign v$G2_13152_out0 = v$RD_6761_out0 && v$RM_12201_out0;
assign v$G2_13156_out0 = v$RD_6765_out0 && v$RM_12205_out0;
assign v$G2_13158_out0 = v$RD_6767_out0 && v$RM_12207_out0;
assign v$G2_13160_out0 = v$RD_6769_out0 && v$RM_12209_out0;
assign v$G2_13163_out0 = v$RD_6772_out0 && v$RM_12212_out0;
assign v$G2_13165_out0 = v$RD_6774_out0 && v$RM_12214_out0;
assign v$G2_13167_out0 = v$RD_6776_out0 && v$RM_12216_out0;
assign v$G2_13169_out0 = v$RD_6778_out0 && v$RM_12218_out0;
assign v$G2_13171_out0 = v$RD_6780_out0 && v$RM_12220_out0;
assign v$G2_13173_out0 = v$RD_6782_out0 && v$RM_12222_out0;
assign v$G2_13175_out0 = v$RD_6784_out0 && v$RM_12224_out0;
assign v$G2_13177_out0 = v$RD_6786_out0 && v$RM_12226_out0;
assign v$G2_13179_out0 = v$RD_6788_out0 && v$RM_12228_out0;
assign v$S_4679_out0 = v$S_9308_out0;
assign v$S_4694_out0 = v$S_9772_out0;
assign v$CARRY_5295_out0 = v$G2_12686_out0;
assign v$CARRY_5297_out0 = v$G2_12688_out0;
assign v$CARRY_5301_out0 = v$G2_12692_out0;
assign v$CARRY_5303_out0 = v$G2_12694_out0;
assign v$CARRY_5305_out0 = v$G2_12696_out0;
assign v$CARRY_5308_out0 = v$G2_12699_out0;
assign v$CARRY_5310_out0 = v$G2_12701_out0;
assign v$CARRY_5312_out0 = v$G2_12703_out0;
assign v$CARRY_5314_out0 = v$G2_12705_out0;
assign v$CARRY_5316_out0 = v$G2_12707_out0;
assign v$CARRY_5318_out0 = v$G2_12709_out0;
assign v$CARRY_5320_out0 = v$G2_12711_out0;
assign v$CARRY_5322_out0 = v$G2_12713_out0;
assign v$CARRY_5324_out0 = v$G2_12715_out0;
assign v$CARRY_5759_out0 = v$G2_13150_out0;
assign v$CARRY_5761_out0 = v$G2_13152_out0;
assign v$CARRY_5765_out0 = v$G2_13156_out0;
assign v$CARRY_5767_out0 = v$G2_13158_out0;
assign v$CARRY_5769_out0 = v$G2_13160_out0;
assign v$CARRY_5772_out0 = v$G2_13163_out0;
assign v$CARRY_5774_out0 = v$G2_13165_out0;
assign v$CARRY_5776_out0 = v$G2_13167_out0;
assign v$CARRY_5778_out0 = v$G2_13169_out0;
assign v$CARRY_5780_out0 = v$G2_13171_out0;
assign v$CARRY_5782_out0 = v$G2_13173_out0;
assign v$CARRY_5784_out0 = v$G2_13175_out0;
assign v$CARRY_5786_out0 = v$G2_13177_out0;
assign v$CARRY_5788_out0 = v$G2_13179_out0;
assign v$S_9296_out0 = v$G1_8150_out0;
assign v$S_9298_out0 = v$G1_8152_out0;
assign v$S_9302_out0 = v$G1_8156_out0;
assign v$S_9304_out0 = v$G1_8158_out0;
assign v$S_9306_out0 = v$G1_8160_out0;
assign v$S_9309_out0 = v$G1_8163_out0;
assign v$S_9311_out0 = v$G1_8165_out0;
assign v$S_9313_out0 = v$G1_8167_out0;
assign v$S_9315_out0 = v$G1_8169_out0;
assign v$S_9317_out0 = v$G1_8171_out0;
assign v$S_9319_out0 = v$G1_8173_out0;
assign v$S_9321_out0 = v$G1_8175_out0;
assign v$S_9323_out0 = v$G1_8177_out0;
assign v$S_9325_out0 = v$G1_8179_out0;
assign v$S_9760_out0 = v$G1_8614_out0;
assign v$S_9762_out0 = v$G1_8616_out0;
assign v$S_9766_out0 = v$G1_8620_out0;
assign v$S_9768_out0 = v$G1_8622_out0;
assign v$S_9770_out0 = v$G1_8624_out0;
assign v$S_9773_out0 = v$G1_8627_out0;
assign v$S_9775_out0 = v$G1_8629_out0;
assign v$S_9777_out0 = v$G1_8631_out0;
assign v$S_9779_out0 = v$G1_8633_out0;
assign v$S_9781_out0 = v$G1_8635_out0;
assign v$S_9783_out0 = v$G1_8637_out0;
assign v$S_9785_out0 = v$G1_8639_out0;
assign v$S_9787_out0 = v$G1_8641_out0;
assign v$S_9789_out0 = v$G1_8643_out0;
assign v$CIN_10025_out0 = v$CARRY_5307_out0;
assign v$CIN_10249_out0 = v$CARRY_5771_out0;
assign v$RD_6313_out0 = v$CIN_10025_out0;
assign v$RD_6777_out0 = v$CIN_10249_out0;
assign v$_10775_out0 = { v$_43_out0,v$S_4679_out0 };
assign v$_10776_out0 = { v$_44_out0,v$S_4694_out0 };
assign v$RM_11736_out0 = v$S_9296_out0;
assign v$RM_11738_out0 = v$S_9298_out0;
assign v$RM_11742_out0 = v$S_9302_out0;
assign v$RM_11744_out0 = v$S_9304_out0;
assign v$RM_11746_out0 = v$S_9306_out0;
assign v$RM_11749_out0 = v$S_9309_out0;
assign v$RM_11751_out0 = v$S_9311_out0;
assign v$RM_11753_out0 = v$S_9313_out0;
assign v$RM_11755_out0 = v$S_9315_out0;
assign v$RM_11757_out0 = v$S_9317_out0;
assign v$RM_11759_out0 = v$S_9319_out0;
assign v$RM_11761_out0 = v$S_9321_out0;
assign v$RM_11763_out0 = v$S_9323_out0;
assign v$RM_11765_out0 = v$S_9325_out0;
assign v$RM_12200_out0 = v$S_9760_out0;
assign v$RM_12202_out0 = v$S_9762_out0;
assign v$RM_12206_out0 = v$S_9766_out0;
assign v$RM_12208_out0 = v$S_9768_out0;
assign v$RM_12210_out0 = v$S_9770_out0;
assign v$RM_12213_out0 = v$S_9773_out0;
assign v$RM_12215_out0 = v$S_9775_out0;
assign v$RM_12217_out0 = v$S_9777_out0;
assign v$RM_12219_out0 = v$S_9779_out0;
assign v$RM_12221_out0 = v$S_9781_out0;
assign v$RM_12223_out0 = v$S_9783_out0;
assign v$RM_12225_out0 = v$S_9785_out0;
assign v$RM_12227_out0 = v$S_9787_out0;
assign v$RM_12229_out0 = v$S_9789_out0;
assign v$G1_8168_out0 = ((v$RD_6313_out0 && !v$RM_11753_out0) || (!v$RD_6313_out0) && v$RM_11753_out0);
assign v$G1_8632_out0 = ((v$RD_6777_out0 && !v$RM_12217_out0) || (!v$RD_6777_out0) && v$RM_12217_out0);
assign v$G2_12704_out0 = v$RD_6313_out0 && v$RM_11753_out0;
assign v$G2_13168_out0 = v$RD_6777_out0 && v$RM_12217_out0;
assign v$CARRY_5313_out0 = v$G2_12704_out0;
assign v$CARRY_5777_out0 = v$G2_13168_out0;
assign v$S_9314_out0 = v$G1_8168_out0;
assign v$S_9778_out0 = v$G1_8632_out0;
assign v$S_1436_out0 = v$S_9314_out0;
assign v$S_1660_out0 = v$S_9778_out0;
assign v$G1_4212_out0 = v$CARRY_5313_out0 || v$CARRY_5312_out0;
assign v$G1_4436_out0 = v$CARRY_5777_out0 || v$CARRY_5776_out0;
assign v$COUT_904_out0 = v$G1_4212_out0;
assign v$COUT_1128_out0 = v$G1_4436_out0;
assign v$CIN_10031_out0 = v$COUT_904_out0;
assign v$CIN_10255_out0 = v$COUT_1128_out0;
assign v$RD_6325_out0 = v$CIN_10031_out0;
assign v$RD_6789_out0 = v$CIN_10255_out0;
assign v$G1_8180_out0 = ((v$RD_6325_out0 && !v$RM_11765_out0) || (!v$RD_6325_out0) && v$RM_11765_out0);
assign v$G1_8644_out0 = ((v$RD_6789_out0 && !v$RM_12229_out0) || (!v$RD_6789_out0) && v$RM_12229_out0);
assign v$G2_12716_out0 = v$RD_6325_out0 && v$RM_11765_out0;
assign v$G2_13180_out0 = v$RD_6789_out0 && v$RM_12229_out0;
assign v$CARRY_5325_out0 = v$G2_12716_out0;
assign v$CARRY_5789_out0 = v$G2_13180_out0;
assign v$S_9326_out0 = v$G1_8180_out0;
assign v$S_9790_out0 = v$G1_8644_out0;
assign v$S_1442_out0 = v$S_9326_out0;
assign v$S_1666_out0 = v$S_9790_out0;
assign v$G1_4218_out0 = v$CARRY_5325_out0 || v$CARRY_5324_out0;
assign v$G1_4442_out0 = v$CARRY_5789_out0 || v$CARRY_5788_out0;
assign v$COUT_910_out0 = v$G1_4218_out0;
assign v$COUT_1134_out0 = v$G1_4442_out0;
assign v$_4796_out0 = { v$S_1436_out0,v$S_1442_out0 };
assign v$_4811_out0 = { v$S_1660_out0,v$S_1666_out0 };
assign v$CIN_10026_out0 = v$COUT_910_out0;
assign v$CIN_10250_out0 = v$COUT_1134_out0;
assign v$RD_6315_out0 = v$CIN_10026_out0;
assign v$RD_6779_out0 = v$CIN_10250_out0;
assign v$G1_8170_out0 = ((v$RD_6315_out0 && !v$RM_11755_out0) || (!v$RD_6315_out0) && v$RM_11755_out0);
assign v$G1_8634_out0 = ((v$RD_6779_out0 && !v$RM_12219_out0) || (!v$RD_6779_out0) && v$RM_12219_out0);
assign v$G2_12706_out0 = v$RD_6315_out0 && v$RM_11755_out0;
assign v$G2_13170_out0 = v$RD_6779_out0 && v$RM_12219_out0;
assign v$CARRY_5315_out0 = v$G2_12706_out0;
assign v$CARRY_5779_out0 = v$G2_13170_out0;
assign v$S_9316_out0 = v$G1_8170_out0;
assign v$S_9780_out0 = v$G1_8634_out0;
assign v$S_1437_out0 = v$S_9316_out0;
assign v$S_1661_out0 = v$S_9780_out0;
assign v$G1_4213_out0 = v$CARRY_5315_out0 || v$CARRY_5314_out0;
assign v$G1_4437_out0 = v$CARRY_5779_out0 || v$CARRY_5778_out0;
assign v$COUT_905_out0 = v$G1_4213_out0;
assign v$COUT_1129_out0 = v$G1_4437_out0;
assign v$_2566_out0 = { v$_4796_out0,v$S_1437_out0 };
assign v$_2581_out0 = { v$_4811_out0,v$S_1661_out0 };
assign v$CIN_10021_out0 = v$COUT_905_out0;
assign v$CIN_10245_out0 = v$COUT_1129_out0;
assign v$RD_6304_out0 = v$CIN_10021_out0;
assign v$RD_6768_out0 = v$CIN_10245_out0;
assign v$G1_8159_out0 = ((v$RD_6304_out0 && !v$RM_11744_out0) || (!v$RD_6304_out0) && v$RM_11744_out0);
assign v$G1_8623_out0 = ((v$RD_6768_out0 && !v$RM_12208_out0) || (!v$RD_6768_out0) && v$RM_12208_out0);
assign v$G2_12695_out0 = v$RD_6304_out0 && v$RM_11744_out0;
assign v$G2_13159_out0 = v$RD_6768_out0 && v$RM_12208_out0;
assign v$CARRY_5304_out0 = v$G2_12695_out0;
assign v$CARRY_5768_out0 = v$G2_13159_out0;
assign v$S_9305_out0 = v$G1_8159_out0;
assign v$S_9769_out0 = v$G1_8623_out0;
assign v$S_1432_out0 = v$S_9305_out0;
assign v$S_1656_out0 = v$S_9769_out0;
assign v$G1_4208_out0 = v$CARRY_5304_out0 || v$CARRY_5303_out0;
assign v$G1_4432_out0 = v$CARRY_5768_out0 || v$CARRY_5767_out0;
assign v$COUT_900_out0 = v$G1_4208_out0;
assign v$COUT_1124_out0 = v$G1_4432_out0;
assign v$_7046_out0 = { v$_2566_out0,v$S_1432_out0 };
assign v$_7061_out0 = { v$_2581_out0,v$S_1656_out0 };
assign v$CIN_10020_out0 = v$COUT_900_out0;
assign v$CIN_10244_out0 = v$COUT_1124_out0;
assign v$RD_6302_out0 = v$CIN_10020_out0;
assign v$RD_6766_out0 = v$CIN_10244_out0;
assign v$G1_8157_out0 = ((v$RD_6302_out0 && !v$RM_11742_out0) || (!v$RD_6302_out0) && v$RM_11742_out0);
assign v$G1_8621_out0 = ((v$RD_6766_out0 && !v$RM_12206_out0) || (!v$RD_6766_out0) && v$RM_12206_out0);
assign v$G2_12693_out0 = v$RD_6302_out0 && v$RM_11742_out0;
assign v$G2_13157_out0 = v$RD_6766_out0 && v$RM_12206_out0;
assign v$CARRY_5302_out0 = v$G2_12693_out0;
assign v$CARRY_5766_out0 = v$G2_13157_out0;
assign v$S_9303_out0 = v$G1_8157_out0;
assign v$S_9767_out0 = v$G1_8621_out0;
assign v$S_1431_out0 = v$S_9303_out0;
assign v$S_1655_out0 = v$S_9767_out0;
assign v$G1_4207_out0 = v$CARRY_5302_out0 || v$CARRY_5301_out0;
assign v$G1_4431_out0 = v$CARRY_5766_out0 || v$CARRY_5765_out0;
assign v$COUT_899_out0 = v$G1_4207_out0;
assign v$COUT_1123_out0 = v$G1_4431_out0;
assign v$_13532_out0 = { v$_7046_out0,v$S_1431_out0 };
assign v$_13547_out0 = { v$_7061_out0,v$S_1655_out0 };
assign v$CIN_10027_out0 = v$COUT_899_out0;
assign v$CIN_10251_out0 = v$COUT_1123_out0;
assign v$RD_6317_out0 = v$CIN_10027_out0;
assign v$RD_6781_out0 = v$CIN_10251_out0;
assign v$G1_8172_out0 = ((v$RD_6317_out0 && !v$RM_11757_out0) || (!v$RD_6317_out0) && v$RM_11757_out0);
assign v$G1_8636_out0 = ((v$RD_6781_out0 && !v$RM_12221_out0) || (!v$RD_6781_out0) && v$RM_12221_out0);
assign v$G2_12708_out0 = v$RD_6317_out0 && v$RM_11757_out0;
assign v$G2_13172_out0 = v$RD_6781_out0 && v$RM_12221_out0;
assign v$CARRY_5317_out0 = v$G2_12708_out0;
assign v$CARRY_5781_out0 = v$G2_13172_out0;
assign v$S_9318_out0 = v$G1_8172_out0;
assign v$S_9782_out0 = v$G1_8636_out0;
assign v$S_1438_out0 = v$S_9318_out0;
assign v$S_1662_out0 = v$S_9782_out0;
assign v$G1_4214_out0 = v$CARRY_5317_out0 || v$CARRY_5316_out0;
assign v$G1_4438_out0 = v$CARRY_5781_out0 || v$CARRY_5780_out0;
assign v$COUT_906_out0 = v$G1_4214_out0;
assign v$COUT_1130_out0 = v$G1_4438_out0;
assign v$_3325_out0 = { v$_13532_out0,v$S_1438_out0 };
assign v$_3340_out0 = { v$_13547_out0,v$S_1662_out0 };
assign v$CIN_10028_out0 = v$COUT_906_out0;
assign v$CIN_10252_out0 = v$COUT_1130_out0;
assign v$RD_6319_out0 = v$CIN_10028_out0;
assign v$RD_6783_out0 = v$CIN_10252_out0;
assign v$G1_8174_out0 = ((v$RD_6319_out0 && !v$RM_11759_out0) || (!v$RD_6319_out0) && v$RM_11759_out0);
assign v$G1_8638_out0 = ((v$RD_6783_out0 && !v$RM_12223_out0) || (!v$RD_6783_out0) && v$RM_12223_out0);
assign v$G2_12710_out0 = v$RD_6319_out0 && v$RM_11759_out0;
assign v$G2_13174_out0 = v$RD_6783_out0 && v$RM_12223_out0;
assign v$CARRY_5319_out0 = v$G2_12710_out0;
assign v$CARRY_5783_out0 = v$G2_13174_out0;
assign v$S_9320_out0 = v$G1_8174_out0;
assign v$S_9784_out0 = v$G1_8638_out0;
assign v$S_1439_out0 = v$S_9320_out0;
assign v$S_1663_out0 = v$S_9784_out0;
assign v$G1_4215_out0 = v$CARRY_5319_out0 || v$CARRY_5318_out0;
assign v$G1_4439_out0 = v$CARRY_5783_out0 || v$CARRY_5782_out0;
assign v$COUT_907_out0 = v$G1_4215_out0;
assign v$COUT_1131_out0 = v$G1_4439_out0;
assign v$_7161_out0 = { v$_3325_out0,v$S_1439_out0 };
assign v$_7176_out0 = { v$_3340_out0,v$S_1663_out0 };
assign v$CIN_10030_out0 = v$COUT_907_out0;
assign v$CIN_10254_out0 = v$COUT_1131_out0;
assign v$RD_6323_out0 = v$CIN_10030_out0;
assign v$RD_6787_out0 = v$CIN_10254_out0;
assign v$G1_8178_out0 = ((v$RD_6323_out0 && !v$RM_11763_out0) || (!v$RD_6323_out0) && v$RM_11763_out0);
assign v$G1_8642_out0 = ((v$RD_6787_out0 && !v$RM_12227_out0) || (!v$RD_6787_out0) && v$RM_12227_out0);
assign v$G2_12714_out0 = v$RD_6323_out0 && v$RM_11763_out0;
assign v$G2_13178_out0 = v$RD_6787_out0 && v$RM_12227_out0;
assign v$CARRY_5323_out0 = v$G2_12714_out0;
assign v$CARRY_5787_out0 = v$G2_13178_out0;
assign v$S_9324_out0 = v$G1_8178_out0;
assign v$S_9788_out0 = v$G1_8642_out0;
assign v$S_1441_out0 = v$S_9324_out0;
assign v$S_1665_out0 = v$S_9788_out0;
assign v$G1_4217_out0 = v$CARRY_5323_out0 || v$CARRY_5322_out0;
assign v$G1_4441_out0 = v$CARRY_5787_out0 || v$CARRY_5786_out0;
assign v$COUT_909_out0 = v$G1_4217_out0;
assign v$COUT_1133_out0 = v$G1_4441_out0;
assign v$_4763_out0 = { v$_7161_out0,v$S_1441_out0 };
assign v$_4778_out0 = { v$_7176_out0,v$S_1665_out0 };
assign v$CIN_10023_out0 = v$COUT_909_out0;
assign v$CIN_10247_out0 = v$COUT_1133_out0;
assign v$RD_6309_out0 = v$CIN_10023_out0;
assign v$RD_6773_out0 = v$CIN_10247_out0;
assign v$G1_8164_out0 = ((v$RD_6309_out0 && !v$RM_11749_out0) || (!v$RD_6309_out0) && v$RM_11749_out0);
assign v$G1_8628_out0 = ((v$RD_6773_out0 && !v$RM_12213_out0) || (!v$RD_6773_out0) && v$RM_12213_out0);
assign v$G2_12700_out0 = v$RD_6309_out0 && v$RM_11749_out0;
assign v$G2_13164_out0 = v$RD_6773_out0 && v$RM_12213_out0;
assign v$CARRY_5309_out0 = v$G2_12700_out0;
assign v$CARRY_5773_out0 = v$G2_13164_out0;
assign v$S_9310_out0 = v$G1_8164_out0;
assign v$S_9774_out0 = v$G1_8628_out0;
assign v$S_1434_out0 = v$S_9310_out0;
assign v$S_1658_out0 = v$S_9774_out0;
assign v$G1_4210_out0 = v$CARRY_5309_out0 || v$CARRY_5308_out0;
assign v$G1_4434_out0 = v$CARRY_5773_out0 || v$CARRY_5772_out0;
assign v$COUT_902_out0 = v$G1_4210_out0;
assign v$COUT_1126_out0 = v$G1_4434_out0;
assign v$_6940_out0 = { v$_4763_out0,v$S_1434_out0 };
assign v$_6955_out0 = { v$_4778_out0,v$S_1658_out0 };
assign v$CIN_10024_out0 = v$COUT_902_out0;
assign v$CIN_10248_out0 = v$COUT_1126_out0;
assign v$RD_6311_out0 = v$CIN_10024_out0;
assign v$RD_6775_out0 = v$CIN_10248_out0;
assign v$G1_8166_out0 = ((v$RD_6311_out0 && !v$RM_11751_out0) || (!v$RD_6311_out0) && v$RM_11751_out0);
assign v$G1_8630_out0 = ((v$RD_6775_out0 && !v$RM_12215_out0) || (!v$RD_6775_out0) && v$RM_12215_out0);
assign v$G2_12702_out0 = v$RD_6311_out0 && v$RM_11751_out0;
assign v$G2_13166_out0 = v$RD_6775_out0 && v$RM_12215_out0;
assign v$CARRY_5311_out0 = v$G2_12702_out0;
assign v$CARRY_5775_out0 = v$G2_13166_out0;
assign v$S_9312_out0 = v$G1_8166_out0;
assign v$S_9776_out0 = v$G1_8630_out0;
assign v$S_1435_out0 = v$S_9312_out0;
assign v$S_1659_out0 = v$S_9776_out0;
assign v$G1_4211_out0 = v$CARRY_5311_out0 || v$CARRY_5310_out0;
assign v$G1_4435_out0 = v$CARRY_5775_out0 || v$CARRY_5774_out0;
assign v$COUT_903_out0 = v$G1_4211_out0;
assign v$COUT_1127_out0 = v$G1_4435_out0;
assign v$_5816_out0 = { v$_6940_out0,v$S_1435_out0 };
assign v$_5831_out0 = { v$_6955_out0,v$S_1659_out0 };
assign v$CIN_10029_out0 = v$COUT_903_out0;
assign v$CIN_10253_out0 = v$COUT_1127_out0;
assign v$RD_6321_out0 = v$CIN_10029_out0;
assign v$RD_6785_out0 = v$CIN_10253_out0;
assign v$G1_8176_out0 = ((v$RD_6321_out0 && !v$RM_11761_out0) || (!v$RD_6321_out0) && v$RM_11761_out0);
assign v$G1_8640_out0 = ((v$RD_6785_out0 && !v$RM_12225_out0) || (!v$RD_6785_out0) && v$RM_12225_out0);
assign v$G2_12712_out0 = v$RD_6321_out0 && v$RM_11761_out0;
assign v$G2_13176_out0 = v$RD_6785_out0 && v$RM_12225_out0;
assign v$CARRY_5321_out0 = v$G2_12712_out0;
assign v$CARRY_5785_out0 = v$G2_13176_out0;
assign v$S_9322_out0 = v$G1_8176_out0;
assign v$S_9786_out0 = v$G1_8640_out0;
assign v$S_1440_out0 = v$S_9322_out0;
assign v$S_1664_out0 = v$S_9786_out0;
assign v$G1_4216_out0 = v$CARRY_5321_out0 || v$CARRY_5320_out0;
assign v$G1_4440_out0 = v$CARRY_5785_out0 || v$CARRY_5784_out0;
assign v$COUT_908_out0 = v$G1_4216_out0;
assign v$COUT_1132_out0 = v$G1_4440_out0;
assign v$_2040_out0 = { v$_5816_out0,v$S_1440_out0 };
assign v$_2055_out0 = { v$_5831_out0,v$S_1664_out0 };
assign v$CIN_10017_out0 = v$COUT_908_out0;
assign v$CIN_10241_out0 = v$COUT_1132_out0;
assign v$RD_6296_out0 = v$CIN_10017_out0;
assign v$RD_6760_out0 = v$CIN_10241_out0;
assign v$G1_8151_out0 = ((v$RD_6296_out0 && !v$RM_11736_out0) || (!v$RD_6296_out0) && v$RM_11736_out0);
assign v$G1_8615_out0 = ((v$RD_6760_out0 && !v$RM_12200_out0) || (!v$RD_6760_out0) && v$RM_12200_out0);
assign v$G2_12687_out0 = v$RD_6296_out0 && v$RM_11736_out0;
assign v$G2_13151_out0 = v$RD_6760_out0 && v$RM_12200_out0;
assign v$CARRY_5296_out0 = v$G2_12687_out0;
assign v$CARRY_5760_out0 = v$G2_13151_out0;
assign v$S_9297_out0 = v$G1_8151_out0;
assign v$S_9761_out0 = v$G1_8615_out0;
assign v$S_1428_out0 = v$S_9297_out0;
assign v$S_1652_out0 = v$S_9761_out0;
assign v$G1_4204_out0 = v$CARRY_5296_out0 || v$CARRY_5295_out0;
assign v$G1_4428_out0 = v$CARRY_5760_out0 || v$CARRY_5759_out0;
assign v$COUT_896_out0 = v$G1_4204_out0;
assign v$COUT_1120_out0 = v$G1_4428_out0;
assign v$_2807_out0 = { v$_2040_out0,v$S_1428_out0 };
assign v$_2822_out0 = { v$_2055_out0,v$S_1652_out0 };
assign v$CIN_10022_out0 = v$COUT_896_out0;
assign v$CIN_10246_out0 = v$COUT_1120_out0;
assign v$RD_6306_out0 = v$CIN_10022_out0;
assign v$RD_6770_out0 = v$CIN_10246_out0;
assign v$G1_8161_out0 = ((v$RD_6306_out0 && !v$RM_11746_out0) || (!v$RD_6306_out0) && v$RM_11746_out0);
assign v$G1_8625_out0 = ((v$RD_6770_out0 && !v$RM_12210_out0) || (!v$RD_6770_out0) && v$RM_12210_out0);
assign v$G2_12697_out0 = v$RD_6306_out0 && v$RM_11746_out0;
assign v$G2_13161_out0 = v$RD_6770_out0 && v$RM_12210_out0;
assign v$CARRY_5306_out0 = v$G2_12697_out0;
assign v$CARRY_5770_out0 = v$G2_13161_out0;
assign v$S_9307_out0 = v$G1_8161_out0;
assign v$S_9771_out0 = v$G1_8625_out0;
assign v$S_1433_out0 = v$S_9307_out0;
assign v$S_1657_out0 = v$S_9771_out0;
assign v$G1_4209_out0 = v$CARRY_5306_out0 || v$CARRY_5305_out0;
assign v$G1_4433_out0 = v$CARRY_5770_out0 || v$CARRY_5769_out0;
assign v$COUT_901_out0 = v$G1_4209_out0;
assign v$COUT_1125_out0 = v$G1_4433_out0;
assign v$_1839_out0 = { v$_2807_out0,v$S_1433_out0 };
assign v$_1854_out0 = { v$_2822_out0,v$S_1657_out0 };
assign v$CIN_10018_out0 = v$COUT_901_out0;
assign v$CIN_10242_out0 = v$COUT_1125_out0;
assign v$RD_6298_out0 = v$CIN_10018_out0;
assign v$RD_6762_out0 = v$CIN_10242_out0;
assign v$G1_8153_out0 = ((v$RD_6298_out0 && !v$RM_11738_out0) || (!v$RD_6298_out0) && v$RM_11738_out0);
assign v$G1_8617_out0 = ((v$RD_6762_out0 && !v$RM_12202_out0) || (!v$RD_6762_out0) && v$RM_12202_out0);
assign v$G2_12689_out0 = v$RD_6298_out0 && v$RM_11738_out0;
assign v$G2_13153_out0 = v$RD_6762_out0 && v$RM_12202_out0;
assign v$CARRY_5298_out0 = v$G2_12689_out0;
assign v$CARRY_5762_out0 = v$G2_13153_out0;
assign v$S_9299_out0 = v$G1_8153_out0;
assign v$S_9763_out0 = v$G1_8617_out0;
assign v$S_1429_out0 = v$S_9299_out0;
assign v$S_1653_out0 = v$S_9763_out0;
assign v$G1_4205_out0 = v$CARRY_5298_out0 || v$CARRY_5297_out0;
assign v$G1_4429_out0 = v$CARRY_5762_out0 || v$CARRY_5761_out0;
assign v$COUT_897_out0 = v$G1_4205_out0;
assign v$COUT_1121_out0 = v$G1_4429_out0;
assign v$_4563_out0 = { v$_1839_out0,v$S_1429_out0 };
assign v$_4578_out0 = { v$_1854_out0,v$S_1653_out0 };
assign v$RM_3566_out0 = v$COUT_897_out0;
assign v$RM_3790_out0 = v$COUT_1121_out0;
assign v$RM_11739_out0 = v$RM_3566_out0;
assign v$RM_12203_out0 = v$RM_3790_out0;
assign v$G1_8154_out0 = ((v$RD_6299_out0 && !v$RM_11739_out0) || (!v$RD_6299_out0) && v$RM_11739_out0);
assign v$G1_8618_out0 = ((v$RD_6763_out0 && !v$RM_12203_out0) || (!v$RD_6763_out0) && v$RM_12203_out0);
assign v$G2_12690_out0 = v$RD_6299_out0 && v$RM_11739_out0;
assign v$G2_13154_out0 = v$RD_6763_out0 && v$RM_12203_out0;
assign v$CARRY_5299_out0 = v$G2_12690_out0;
assign v$CARRY_5763_out0 = v$G2_13154_out0;
assign v$S_9300_out0 = v$G1_8154_out0;
assign v$S_9764_out0 = v$G1_8618_out0;
assign v$RM_11740_out0 = v$S_9300_out0;
assign v$RM_12204_out0 = v$S_9764_out0;
assign v$G1_8155_out0 = ((v$RD_6300_out0 && !v$RM_11740_out0) || (!v$RD_6300_out0) && v$RM_11740_out0);
assign v$G1_8619_out0 = ((v$RD_6764_out0 && !v$RM_12204_out0) || (!v$RD_6764_out0) && v$RM_12204_out0);
assign v$G2_12691_out0 = v$RD_6300_out0 && v$RM_11740_out0;
assign v$G2_13155_out0 = v$RD_6764_out0 && v$RM_12204_out0;
assign v$CARRY_5300_out0 = v$G2_12691_out0;
assign v$CARRY_5764_out0 = v$G2_13155_out0;
assign v$S_9301_out0 = v$G1_8155_out0;
assign v$S_9765_out0 = v$G1_8619_out0;
assign v$S_1430_out0 = v$S_9301_out0;
assign v$S_1654_out0 = v$S_9765_out0;
assign v$G1_4206_out0 = v$CARRY_5300_out0 || v$CARRY_5299_out0;
assign v$G1_4430_out0 = v$CARRY_5764_out0 || v$CARRY_5763_out0;
assign v$COUT_898_out0 = v$G1_4206_out0;
assign v$COUT_1122_out0 = v$G1_4430_out0;
assign v$_10665_out0 = { v$_4563_out0,v$S_1430_out0 };
assign v$_10680_out0 = { v$_4578_out0,v$S_1654_out0 };
assign v$_10960_out0 = { v$_10665_out0,v$COUT_898_out0 };
assign v$_10975_out0 = { v$_10680_out0,v$COUT_1122_out0 };
assign v$COUT_10930_out0 = v$_10960_out0;
assign v$COUT_10945_out0 = v$_10975_out0;
assign v$CIN_2360_out0 = v$COUT_10930_out0;
assign v$CIN_2375_out0 = v$COUT_10945_out0;
assign v$_473_out0 = v$CIN_2360_out0[8:8];
assign v$_488_out0 = v$CIN_2375_out0[8:8];
assign v$_1778_out0 = v$CIN_2360_out0[6:6];
assign v$_1793_out0 = v$CIN_2375_out0[6:6];
assign v$_2160_out0 = v$CIN_2360_out0[3:3];
assign v$_2175_out0 = v$CIN_2375_out0[3:3];
assign v$_2199_out0 = v$CIN_2360_out0[15:15];
assign v$_2213_out0 = v$CIN_2375_out0[15:15];
assign v$_2507_out0 = v$CIN_2360_out0[0:0];
assign v$_2522_out0 = v$CIN_2375_out0[0:0];
assign v$_3056_out0 = v$CIN_2360_out0[9:9];
assign v$_3071_out0 = v$CIN_2375_out0[9:9];
assign v$_3090_out0 = v$CIN_2360_out0[2:2];
assign v$_3105_out0 = v$CIN_2375_out0[2:2];
assign v$_3144_out0 = v$CIN_2360_out0[7:7];
assign v$_3159_out0 = v$CIN_2375_out0[7:7];
assign v$_3828_out0 = v$CIN_2360_out0[1:1];
assign v$_3843_out0 = v$CIN_2375_out0[1:1];
assign v$_3866_out0 = v$CIN_2360_out0[10:10];
assign v$_3881_out0 = v$CIN_2375_out0[10:10];
assign v$_6805_out0 = v$CIN_2360_out0[11:11];
assign v$_6820_out0 = v$CIN_2375_out0[11:11];
assign v$_7649_out0 = v$CIN_2360_out0[12:12];
assign v$_7664_out0 = v$CIN_2375_out0[12:12];
assign v$_8704_out0 = v$CIN_2360_out0[13:13];
assign v$_8719_out0 = v$CIN_2375_out0[13:13];
assign v$_8774_out0 = v$CIN_2360_out0[14:14];
assign v$_8789_out0 = v$CIN_2375_out0[14:14];
assign v$_10724_out0 = v$CIN_2360_out0[5:5];
assign v$_10739_out0 = v$CIN_2375_out0[5:5];
assign v$_13453_out0 = v$CIN_2360_out0[4:4];
assign v$_13468_out0 = v$CIN_2375_out0[4:4];
assign v$RM_3429_out0 = v$_7649_out0;
assign v$RM_3430_out0 = v$_8774_out0;
assign v$RM_3432_out0 = v$_10724_out0;
assign v$RM_3433_out0 = v$_13453_out0;
assign v$RM_3434_out0 = v$_8704_out0;
assign v$RM_3435_out0 = v$_3056_out0;
assign v$RM_3436_out0 = v$_3866_out0;
assign v$RM_3437_out0 = v$_3828_out0;
assign v$RM_3438_out0 = v$_2160_out0;
assign v$RM_3439_out0 = v$_1778_out0;
assign v$RM_3440_out0 = v$_3144_out0;
assign v$RM_3441_out0 = v$_6805_out0;
assign v$RM_3442_out0 = v$_473_out0;
assign v$RM_3443_out0 = v$_3090_out0;
assign v$RM_3653_out0 = v$_7664_out0;
assign v$RM_3654_out0 = v$_8789_out0;
assign v$RM_3656_out0 = v$_10739_out0;
assign v$RM_3657_out0 = v$_13468_out0;
assign v$RM_3658_out0 = v$_8719_out0;
assign v$RM_3659_out0 = v$_3071_out0;
assign v$RM_3660_out0 = v$_3881_out0;
assign v$RM_3661_out0 = v$_3843_out0;
assign v$RM_3662_out0 = v$_2175_out0;
assign v$RM_3663_out0 = v$_1793_out0;
assign v$RM_3664_out0 = v$_3159_out0;
assign v$RM_3665_out0 = v$_6820_out0;
assign v$RM_3666_out0 = v$_488_out0;
assign v$RM_3667_out0 = v$_3105_out0;
assign v$CIN_9884_out0 = v$_2199_out0;
assign v$CIN_10108_out0 = v$_2213_out0;
assign v$RM_11468_out0 = v$_2507_out0;
assign v$RM_11932_out0 = v$_2522_out0;
assign v$RD_6021_out0 = v$CIN_9884_out0;
assign v$RD_6485_out0 = v$CIN_10108_out0;
assign v$G1_7883_out0 = ((v$RD_6028_out0 && !v$RM_11468_out0) || (!v$RD_6028_out0) && v$RM_11468_out0);
assign v$G1_8347_out0 = ((v$RD_6492_out0 && !v$RM_11932_out0) || (!v$RD_6492_out0) && v$RM_11932_out0);
assign v$RM_11456_out0 = v$RM_3429_out0;
assign v$RM_11458_out0 = v$RM_3430_out0;
assign v$RM_11462_out0 = v$RM_3432_out0;
assign v$RM_11464_out0 = v$RM_3433_out0;
assign v$RM_11466_out0 = v$RM_3434_out0;
assign v$RM_11469_out0 = v$RM_3435_out0;
assign v$RM_11471_out0 = v$RM_3436_out0;
assign v$RM_11473_out0 = v$RM_3437_out0;
assign v$RM_11475_out0 = v$RM_3438_out0;
assign v$RM_11477_out0 = v$RM_3439_out0;
assign v$RM_11479_out0 = v$RM_3440_out0;
assign v$RM_11481_out0 = v$RM_3441_out0;
assign v$RM_11483_out0 = v$RM_3442_out0;
assign v$RM_11485_out0 = v$RM_3443_out0;
assign v$RM_11920_out0 = v$RM_3653_out0;
assign v$RM_11922_out0 = v$RM_3654_out0;
assign v$RM_11926_out0 = v$RM_3656_out0;
assign v$RM_11928_out0 = v$RM_3657_out0;
assign v$RM_11930_out0 = v$RM_3658_out0;
assign v$RM_11933_out0 = v$RM_3659_out0;
assign v$RM_11935_out0 = v$RM_3660_out0;
assign v$RM_11937_out0 = v$RM_3661_out0;
assign v$RM_11939_out0 = v$RM_3662_out0;
assign v$RM_11941_out0 = v$RM_3663_out0;
assign v$RM_11943_out0 = v$RM_3664_out0;
assign v$RM_11945_out0 = v$RM_3665_out0;
assign v$RM_11947_out0 = v$RM_3666_out0;
assign v$RM_11949_out0 = v$RM_3667_out0;
assign v$G2_12419_out0 = v$RD_6028_out0 && v$RM_11468_out0;
assign v$G2_12883_out0 = v$RD_6492_out0 && v$RM_11932_out0;
assign v$CARRY_5028_out0 = v$G2_12419_out0;
assign v$CARRY_5492_out0 = v$G2_12883_out0;
assign v$G1_7871_out0 = ((v$RD_6016_out0 && !v$RM_11456_out0) || (!v$RD_6016_out0) && v$RM_11456_out0);
assign v$G1_7873_out0 = ((v$RD_6018_out0 && !v$RM_11458_out0) || (!v$RD_6018_out0) && v$RM_11458_out0);
assign v$G1_7877_out0 = ((v$RD_6022_out0 && !v$RM_11462_out0) || (!v$RD_6022_out0) && v$RM_11462_out0);
assign v$G1_7879_out0 = ((v$RD_6024_out0 && !v$RM_11464_out0) || (!v$RD_6024_out0) && v$RM_11464_out0);
assign v$G1_7881_out0 = ((v$RD_6026_out0 && !v$RM_11466_out0) || (!v$RD_6026_out0) && v$RM_11466_out0);
assign v$G1_7884_out0 = ((v$RD_6029_out0 && !v$RM_11469_out0) || (!v$RD_6029_out0) && v$RM_11469_out0);
assign v$G1_7886_out0 = ((v$RD_6031_out0 && !v$RM_11471_out0) || (!v$RD_6031_out0) && v$RM_11471_out0);
assign v$G1_7888_out0 = ((v$RD_6033_out0 && !v$RM_11473_out0) || (!v$RD_6033_out0) && v$RM_11473_out0);
assign v$G1_7890_out0 = ((v$RD_6035_out0 && !v$RM_11475_out0) || (!v$RD_6035_out0) && v$RM_11475_out0);
assign v$G1_7892_out0 = ((v$RD_6037_out0 && !v$RM_11477_out0) || (!v$RD_6037_out0) && v$RM_11477_out0);
assign v$G1_7894_out0 = ((v$RD_6039_out0 && !v$RM_11479_out0) || (!v$RD_6039_out0) && v$RM_11479_out0);
assign v$G1_7896_out0 = ((v$RD_6041_out0 && !v$RM_11481_out0) || (!v$RD_6041_out0) && v$RM_11481_out0);
assign v$G1_7898_out0 = ((v$RD_6043_out0 && !v$RM_11483_out0) || (!v$RD_6043_out0) && v$RM_11483_out0);
assign v$G1_7900_out0 = ((v$RD_6045_out0 && !v$RM_11485_out0) || (!v$RD_6045_out0) && v$RM_11485_out0);
assign v$G1_8335_out0 = ((v$RD_6480_out0 && !v$RM_11920_out0) || (!v$RD_6480_out0) && v$RM_11920_out0);
assign v$G1_8337_out0 = ((v$RD_6482_out0 && !v$RM_11922_out0) || (!v$RD_6482_out0) && v$RM_11922_out0);
assign v$G1_8341_out0 = ((v$RD_6486_out0 && !v$RM_11926_out0) || (!v$RD_6486_out0) && v$RM_11926_out0);
assign v$G1_8343_out0 = ((v$RD_6488_out0 && !v$RM_11928_out0) || (!v$RD_6488_out0) && v$RM_11928_out0);
assign v$G1_8345_out0 = ((v$RD_6490_out0 && !v$RM_11930_out0) || (!v$RD_6490_out0) && v$RM_11930_out0);
assign v$G1_8348_out0 = ((v$RD_6493_out0 && !v$RM_11933_out0) || (!v$RD_6493_out0) && v$RM_11933_out0);
assign v$G1_8350_out0 = ((v$RD_6495_out0 && !v$RM_11935_out0) || (!v$RD_6495_out0) && v$RM_11935_out0);
assign v$G1_8352_out0 = ((v$RD_6497_out0 && !v$RM_11937_out0) || (!v$RD_6497_out0) && v$RM_11937_out0);
assign v$G1_8354_out0 = ((v$RD_6499_out0 && !v$RM_11939_out0) || (!v$RD_6499_out0) && v$RM_11939_out0);
assign v$G1_8356_out0 = ((v$RD_6501_out0 && !v$RM_11941_out0) || (!v$RD_6501_out0) && v$RM_11941_out0);
assign v$G1_8358_out0 = ((v$RD_6503_out0 && !v$RM_11943_out0) || (!v$RD_6503_out0) && v$RM_11943_out0);
assign v$G1_8360_out0 = ((v$RD_6505_out0 && !v$RM_11945_out0) || (!v$RD_6505_out0) && v$RM_11945_out0);
assign v$G1_8362_out0 = ((v$RD_6507_out0 && !v$RM_11947_out0) || (!v$RD_6507_out0) && v$RM_11947_out0);
assign v$G1_8364_out0 = ((v$RD_6509_out0 && !v$RM_11949_out0) || (!v$RD_6509_out0) && v$RM_11949_out0);
assign v$S_9029_out0 = v$G1_7883_out0;
assign v$S_9493_out0 = v$G1_8347_out0;
assign v$G2_12407_out0 = v$RD_6016_out0 && v$RM_11456_out0;
assign v$G2_12409_out0 = v$RD_6018_out0 && v$RM_11458_out0;
assign v$G2_12413_out0 = v$RD_6022_out0 && v$RM_11462_out0;
assign v$G2_12415_out0 = v$RD_6024_out0 && v$RM_11464_out0;
assign v$G2_12417_out0 = v$RD_6026_out0 && v$RM_11466_out0;
assign v$G2_12420_out0 = v$RD_6029_out0 && v$RM_11469_out0;
assign v$G2_12422_out0 = v$RD_6031_out0 && v$RM_11471_out0;
assign v$G2_12424_out0 = v$RD_6033_out0 && v$RM_11473_out0;
assign v$G2_12426_out0 = v$RD_6035_out0 && v$RM_11475_out0;
assign v$G2_12428_out0 = v$RD_6037_out0 && v$RM_11477_out0;
assign v$G2_12430_out0 = v$RD_6039_out0 && v$RM_11479_out0;
assign v$G2_12432_out0 = v$RD_6041_out0 && v$RM_11481_out0;
assign v$G2_12434_out0 = v$RD_6043_out0 && v$RM_11483_out0;
assign v$G2_12436_out0 = v$RD_6045_out0 && v$RM_11485_out0;
assign v$G2_12871_out0 = v$RD_6480_out0 && v$RM_11920_out0;
assign v$G2_12873_out0 = v$RD_6482_out0 && v$RM_11922_out0;
assign v$G2_12877_out0 = v$RD_6486_out0 && v$RM_11926_out0;
assign v$G2_12879_out0 = v$RD_6488_out0 && v$RM_11928_out0;
assign v$G2_12881_out0 = v$RD_6490_out0 && v$RM_11930_out0;
assign v$G2_12884_out0 = v$RD_6493_out0 && v$RM_11933_out0;
assign v$G2_12886_out0 = v$RD_6495_out0 && v$RM_11935_out0;
assign v$G2_12888_out0 = v$RD_6497_out0 && v$RM_11937_out0;
assign v$G2_12890_out0 = v$RD_6499_out0 && v$RM_11939_out0;
assign v$G2_12892_out0 = v$RD_6501_out0 && v$RM_11941_out0;
assign v$G2_12894_out0 = v$RD_6503_out0 && v$RM_11943_out0;
assign v$G2_12896_out0 = v$RD_6505_out0 && v$RM_11945_out0;
assign v$G2_12898_out0 = v$RD_6507_out0 && v$RM_11947_out0;
assign v$G2_12900_out0 = v$RD_6509_out0 && v$RM_11949_out0;
assign v$S_4670_out0 = v$S_9029_out0;
assign v$S_4685_out0 = v$S_9493_out0;
assign v$CARRY_5016_out0 = v$G2_12407_out0;
assign v$CARRY_5018_out0 = v$G2_12409_out0;
assign v$CARRY_5022_out0 = v$G2_12413_out0;
assign v$CARRY_5024_out0 = v$G2_12415_out0;
assign v$CARRY_5026_out0 = v$G2_12417_out0;
assign v$CARRY_5029_out0 = v$G2_12420_out0;
assign v$CARRY_5031_out0 = v$G2_12422_out0;
assign v$CARRY_5033_out0 = v$G2_12424_out0;
assign v$CARRY_5035_out0 = v$G2_12426_out0;
assign v$CARRY_5037_out0 = v$G2_12428_out0;
assign v$CARRY_5039_out0 = v$G2_12430_out0;
assign v$CARRY_5041_out0 = v$G2_12432_out0;
assign v$CARRY_5043_out0 = v$G2_12434_out0;
assign v$CARRY_5045_out0 = v$G2_12436_out0;
assign v$CARRY_5480_out0 = v$G2_12871_out0;
assign v$CARRY_5482_out0 = v$G2_12873_out0;
assign v$CARRY_5486_out0 = v$G2_12877_out0;
assign v$CARRY_5488_out0 = v$G2_12879_out0;
assign v$CARRY_5490_out0 = v$G2_12881_out0;
assign v$CARRY_5493_out0 = v$G2_12884_out0;
assign v$CARRY_5495_out0 = v$G2_12886_out0;
assign v$CARRY_5497_out0 = v$G2_12888_out0;
assign v$CARRY_5499_out0 = v$G2_12890_out0;
assign v$CARRY_5501_out0 = v$G2_12892_out0;
assign v$CARRY_5503_out0 = v$G2_12894_out0;
assign v$CARRY_5505_out0 = v$G2_12896_out0;
assign v$CARRY_5507_out0 = v$G2_12898_out0;
assign v$CARRY_5509_out0 = v$G2_12900_out0;
assign v$S_9017_out0 = v$G1_7871_out0;
assign v$S_9019_out0 = v$G1_7873_out0;
assign v$S_9023_out0 = v$G1_7877_out0;
assign v$S_9025_out0 = v$G1_7879_out0;
assign v$S_9027_out0 = v$G1_7881_out0;
assign v$S_9030_out0 = v$G1_7884_out0;
assign v$S_9032_out0 = v$G1_7886_out0;
assign v$S_9034_out0 = v$G1_7888_out0;
assign v$S_9036_out0 = v$G1_7890_out0;
assign v$S_9038_out0 = v$G1_7892_out0;
assign v$S_9040_out0 = v$G1_7894_out0;
assign v$S_9042_out0 = v$G1_7896_out0;
assign v$S_9044_out0 = v$G1_7898_out0;
assign v$S_9046_out0 = v$G1_7900_out0;
assign v$S_9481_out0 = v$G1_8335_out0;
assign v$S_9483_out0 = v$G1_8337_out0;
assign v$S_9487_out0 = v$G1_8341_out0;
assign v$S_9489_out0 = v$G1_8343_out0;
assign v$S_9491_out0 = v$G1_8345_out0;
assign v$S_9494_out0 = v$G1_8348_out0;
assign v$S_9496_out0 = v$G1_8350_out0;
assign v$S_9498_out0 = v$G1_8352_out0;
assign v$S_9500_out0 = v$G1_8354_out0;
assign v$S_9502_out0 = v$G1_8356_out0;
assign v$S_9504_out0 = v$G1_8358_out0;
assign v$S_9506_out0 = v$G1_8360_out0;
assign v$S_9508_out0 = v$G1_8362_out0;
assign v$S_9510_out0 = v$G1_8364_out0;
assign v$CIN_9890_out0 = v$CARRY_5028_out0;
assign v$CIN_10114_out0 = v$CARRY_5492_out0;
assign v$_2191_out0 = { v$_10775_out0,v$S_4670_out0 };
assign v$_2192_out0 = { v$_10776_out0,v$S_4685_out0 };
assign v$RD_6034_out0 = v$CIN_9890_out0;
assign v$RD_6498_out0 = v$CIN_10114_out0;
assign v$RM_11457_out0 = v$S_9017_out0;
assign v$RM_11459_out0 = v$S_9019_out0;
assign v$RM_11463_out0 = v$S_9023_out0;
assign v$RM_11465_out0 = v$S_9025_out0;
assign v$RM_11467_out0 = v$S_9027_out0;
assign v$RM_11470_out0 = v$S_9030_out0;
assign v$RM_11472_out0 = v$S_9032_out0;
assign v$RM_11474_out0 = v$S_9034_out0;
assign v$RM_11476_out0 = v$S_9036_out0;
assign v$RM_11478_out0 = v$S_9038_out0;
assign v$RM_11480_out0 = v$S_9040_out0;
assign v$RM_11482_out0 = v$S_9042_out0;
assign v$RM_11484_out0 = v$S_9044_out0;
assign v$RM_11486_out0 = v$S_9046_out0;
assign v$RM_11921_out0 = v$S_9481_out0;
assign v$RM_11923_out0 = v$S_9483_out0;
assign v$RM_11927_out0 = v$S_9487_out0;
assign v$RM_11929_out0 = v$S_9489_out0;
assign v$RM_11931_out0 = v$S_9491_out0;
assign v$RM_11934_out0 = v$S_9494_out0;
assign v$RM_11936_out0 = v$S_9496_out0;
assign v$RM_11938_out0 = v$S_9498_out0;
assign v$RM_11940_out0 = v$S_9500_out0;
assign v$RM_11942_out0 = v$S_9502_out0;
assign v$RM_11944_out0 = v$S_9504_out0;
assign v$RM_11946_out0 = v$S_9506_out0;
assign v$RM_11948_out0 = v$S_9508_out0;
assign v$RM_11950_out0 = v$S_9510_out0;
assign v$G1_7889_out0 = ((v$RD_6034_out0 && !v$RM_11474_out0) || (!v$RD_6034_out0) && v$RM_11474_out0);
assign v$G1_8353_out0 = ((v$RD_6498_out0 && !v$RM_11938_out0) || (!v$RD_6498_out0) && v$RM_11938_out0);
assign v$G2_12425_out0 = v$RD_6034_out0 && v$RM_11474_out0;
assign v$G2_12889_out0 = v$RD_6498_out0 && v$RM_11938_out0;
assign v$CARRY_5034_out0 = v$G2_12425_out0;
assign v$CARRY_5498_out0 = v$G2_12889_out0;
assign v$S_9035_out0 = v$G1_7889_out0;
assign v$S_9499_out0 = v$G1_8353_out0;
assign v$S_1301_out0 = v$S_9035_out0;
assign v$S_1525_out0 = v$S_9499_out0;
assign v$G1_4077_out0 = v$CARRY_5034_out0 || v$CARRY_5033_out0;
assign v$G1_4301_out0 = v$CARRY_5498_out0 || v$CARRY_5497_out0;
assign v$COUT_769_out0 = v$G1_4077_out0;
assign v$COUT_993_out0 = v$G1_4301_out0;
assign v$CIN_9896_out0 = v$COUT_769_out0;
assign v$CIN_10120_out0 = v$COUT_993_out0;
assign v$RD_6046_out0 = v$CIN_9896_out0;
assign v$RD_6510_out0 = v$CIN_10120_out0;
assign v$G1_7901_out0 = ((v$RD_6046_out0 && !v$RM_11486_out0) || (!v$RD_6046_out0) && v$RM_11486_out0);
assign v$G1_8365_out0 = ((v$RD_6510_out0 && !v$RM_11950_out0) || (!v$RD_6510_out0) && v$RM_11950_out0);
assign v$G2_12437_out0 = v$RD_6046_out0 && v$RM_11486_out0;
assign v$G2_12901_out0 = v$RD_6510_out0 && v$RM_11950_out0;
assign v$CARRY_5046_out0 = v$G2_12437_out0;
assign v$CARRY_5510_out0 = v$G2_12901_out0;
assign v$S_9047_out0 = v$G1_7901_out0;
assign v$S_9511_out0 = v$G1_8365_out0;
assign v$S_1307_out0 = v$S_9047_out0;
assign v$S_1531_out0 = v$S_9511_out0;
assign v$G1_4083_out0 = v$CARRY_5046_out0 || v$CARRY_5045_out0;
assign v$G1_4307_out0 = v$CARRY_5510_out0 || v$CARRY_5509_out0;
assign v$COUT_775_out0 = v$G1_4083_out0;
assign v$COUT_999_out0 = v$G1_4307_out0;
assign v$_4787_out0 = { v$S_1301_out0,v$S_1307_out0 };
assign v$_4802_out0 = { v$S_1525_out0,v$S_1531_out0 };
assign v$CIN_9891_out0 = v$COUT_775_out0;
assign v$CIN_10115_out0 = v$COUT_999_out0;
assign v$RD_6036_out0 = v$CIN_9891_out0;
assign v$RD_6500_out0 = v$CIN_10115_out0;
assign v$G1_7891_out0 = ((v$RD_6036_out0 && !v$RM_11476_out0) || (!v$RD_6036_out0) && v$RM_11476_out0);
assign v$G1_8355_out0 = ((v$RD_6500_out0 && !v$RM_11940_out0) || (!v$RD_6500_out0) && v$RM_11940_out0);
assign v$G2_12427_out0 = v$RD_6036_out0 && v$RM_11476_out0;
assign v$G2_12891_out0 = v$RD_6500_out0 && v$RM_11940_out0;
assign v$CARRY_5036_out0 = v$G2_12427_out0;
assign v$CARRY_5500_out0 = v$G2_12891_out0;
assign v$S_9037_out0 = v$G1_7891_out0;
assign v$S_9501_out0 = v$G1_8355_out0;
assign v$S_1302_out0 = v$S_9037_out0;
assign v$S_1526_out0 = v$S_9501_out0;
assign v$G1_4078_out0 = v$CARRY_5036_out0 || v$CARRY_5035_out0;
assign v$G1_4302_out0 = v$CARRY_5500_out0 || v$CARRY_5499_out0;
assign v$COUT_770_out0 = v$G1_4078_out0;
assign v$COUT_994_out0 = v$G1_4302_out0;
assign v$_2557_out0 = { v$_4787_out0,v$S_1302_out0 };
assign v$_2572_out0 = { v$_4802_out0,v$S_1526_out0 };
assign v$CIN_9886_out0 = v$COUT_770_out0;
assign v$CIN_10110_out0 = v$COUT_994_out0;
assign v$RD_6025_out0 = v$CIN_9886_out0;
assign v$RD_6489_out0 = v$CIN_10110_out0;
assign v$G1_7880_out0 = ((v$RD_6025_out0 && !v$RM_11465_out0) || (!v$RD_6025_out0) && v$RM_11465_out0);
assign v$G1_8344_out0 = ((v$RD_6489_out0 && !v$RM_11929_out0) || (!v$RD_6489_out0) && v$RM_11929_out0);
assign v$G2_12416_out0 = v$RD_6025_out0 && v$RM_11465_out0;
assign v$G2_12880_out0 = v$RD_6489_out0 && v$RM_11929_out0;
assign v$CARRY_5025_out0 = v$G2_12416_out0;
assign v$CARRY_5489_out0 = v$G2_12880_out0;
assign v$S_9026_out0 = v$G1_7880_out0;
assign v$S_9490_out0 = v$G1_8344_out0;
assign v$S_1297_out0 = v$S_9026_out0;
assign v$S_1521_out0 = v$S_9490_out0;
assign v$G1_4073_out0 = v$CARRY_5025_out0 || v$CARRY_5024_out0;
assign v$G1_4297_out0 = v$CARRY_5489_out0 || v$CARRY_5488_out0;
assign v$COUT_765_out0 = v$G1_4073_out0;
assign v$COUT_989_out0 = v$G1_4297_out0;
assign v$_7037_out0 = { v$_2557_out0,v$S_1297_out0 };
assign v$_7052_out0 = { v$_2572_out0,v$S_1521_out0 };
assign v$CIN_9885_out0 = v$COUT_765_out0;
assign v$CIN_10109_out0 = v$COUT_989_out0;
assign v$RD_6023_out0 = v$CIN_9885_out0;
assign v$RD_6487_out0 = v$CIN_10109_out0;
assign v$G1_7878_out0 = ((v$RD_6023_out0 && !v$RM_11463_out0) || (!v$RD_6023_out0) && v$RM_11463_out0);
assign v$G1_8342_out0 = ((v$RD_6487_out0 && !v$RM_11927_out0) || (!v$RD_6487_out0) && v$RM_11927_out0);
assign v$G2_12414_out0 = v$RD_6023_out0 && v$RM_11463_out0;
assign v$G2_12878_out0 = v$RD_6487_out0 && v$RM_11927_out0;
assign v$CARRY_5023_out0 = v$G2_12414_out0;
assign v$CARRY_5487_out0 = v$G2_12878_out0;
assign v$S_9024_out0 = v$G1_7878_out0;
assign v$S_9488_out0 = v$G1_8342_out0;
assign v$S_1296_out0 = v$S_9024_out0;
assign v$S_1520_out0 = v$S_9488_out0;
assign v$G1_4072_out0 = v$CARRY_5023_out0 || v$CARRY_5022_out0;
assign v$G1_4296_out0 = v$CARRY_5487_out0 || v$CARRY_5486_out0;
assign v$COUT_764_out0 = v$G1_4072_out0;
assign v$COUT_988_out0 = v$G1_4296_out0;
assign v$_13523_out0 = { v$_7037_out0,v$S_1296_out0 };
assign v$_13538_out0 = { v$_7052_out0,v$S_1520_out0 };
assign v$CIN_9892_out0 = v$COUT_764_out0;
assign v$CIN_10116_out0 = v$COUT_988_out0;
assign v$RD_6038_out0 = v$CIN_9892_out0;
assign v$RD_6502_out0 = v$CIN_10116_out0;
assign v$G1_7893_out0 = ((v$RD_6038_out0 && !v$RM_11478_out0) || (!v$RD_6038_out0) && v$RM_11478_out0);
assign v$G1_8357_out0 = ((v$RD_6502_out0 && !v$RM_11942_out0) || (!v$RD_6502_out0) && v$RM_11942_out0);
assign v$G2_12429_out0 = v$RD_6038_out0 && v$RM_11478_out0;
assign v$G2_12893_out0 = v$RD_6502_out0 && v$RM_11942_out0;
assign v$CARRY_5038_out0 = v$G2_12429_out0;
assign v$CARRY_5502_out0 = v$G2_12893_out0;
assign v$S_9039_out0 = v$G1_7893_out0;
assign v$S_9503_out0 = v$G1_8357_out0;
assign v$S_1303_out0 = v$S_9039_out0;
assign v$S_1527_out0 = v$S_9503_out0;
assign v$G1_4079_out0 = v$CARRY_5038_out0 || v$CARRY_5037_out0;
assign v$G1_4303_out0 = v$CARRY_5502_out0 || v$CARRY_5501_out0;
assign v$COUT_771_out0 = v$G1_4079_out0;
assign v$COUT_995_out0 = v$G1_4303_out0;
assign v$_3316_out0 = { v$_13523_out0,v$S_1303_out0 };
assign v$_3331_out0 = { v$_13538_out0,v$S_1527_out0 };
assign v$CIN_9893_out0 = v$COUT_771_out0;
assign v$CIN_10117_out0 = v$COUT_995_out0;
assign v$RD_6040_out0 = v$CIN_9893_out0;
assign v$RD_6504_out0 = v$CIN_10117_out0;
assign v$G1_7895_out0 = ((v$RD_6040_out0 && !v$RM_11480_out0) || (!v$RD_6040_out0) && v$RM_11480_out0);
assign v$G1_8359_out0 = ((v$RD_6504_out0 && !v$RM_11944_out0) || (!v$RD_6504_out0) && v$RM_11944_out0);
assign v$G2_12431_out0 = v$RD_6040_out0 && v$RM_11480_out0;
assign v$G2_12895_out0 = v$RD_6504_out0 && v$RM_11944_out0;
assign v$CARRY_5040_out0 = v$G2_12431_out0;
assign v$CARRY_5504_out0 = v$G2_12895_out0;
assign v$S_9041_out0 = v$G1_7895_out0;
assign v$S_9505_out0 = v$G1_8359_out0;
assign v$S_1304_out0 = v$S_9041_out0;
assign v$S_1528_out0 = v$S_9505_out0;
assign v$G1_4080_out0 = v$CARRY_5040_out0 || v$CARRY_5039_out0;
assign v$G1_4304_out0 = v$CARRY_5504_out0 || v$CARRY_5503_out0;
assign v$COUT_772_out0 = v$G1_4080_out0;
assign v$COUT_996_out0 = v$G1_4304_out0;
assign v$_7152_out0 = { v$_3316_out0,v$S_1304_out0 };
assign v$_7167_out0 = { v$_3331_out0,v$S_1528_out0 };
assign v$CIN_9895_out0 = v$COUT_772_out0;
assign v$CIN_10119_out0 = v$COUT_996_out0;
assign v$RD_6044_out0 = v$CIN_9895_out0;
assign v$RD_6508_out0 = v$CIN_10119_out0;
assign v$G1_7899_out0 = ((v$RD_6044_out0 && !v$RM_11484_out0) || (!v$RD_6044_out0) && v$RM_11484_out0);
assign v$G1_8363_out0 = ((v$RD_6508_out0 && !v$RM_11948_out0) || (!v$RD_6508_out0) && v$RM_11948_out0);
assign v$G2_12435_out0 = v$RD_6044_out0 && v$RM_11484_out0;
assign v$G2_12899_out0 = v$RD_6508_out0 && v$RM_11948_out0;
assign v$CARRY_5044_out0 = v$G2_12435_out0;
assign v$CARRY_5508_out0 = v$G2_12899_out0;
assign v$S_9045_out0 = v$G1_7899_out0;
assign v$S_9509_out0 = v$G1_8363_out0;
assign v$S_1306_out0 = v$S_9045_out0;
assign v$S_1530_out0 = v$S_9509_out0;
assign v$G1_4082_out0 = v$CARRY_5044_out0 || v$CARRY_5043_out0;
assign v$G1_4306_out0 = v$CARRY_5508_out0 || v$CARRY_5507_out0;
assign v$COUT_774_out0 = v$G1_4082_out0;
assign v$COUT_998_out0 = v$G1_4306_out0;
assign v$_4754_out0 = { v$_7152_out0,v$S_1306_out0 };
assign v$_4769_out0 = { v$_7167_out0,v$S_1530_out0 };
assign v$CIN_9888_out0 = v$COUT_774_out0;
assign v$CIN_10112_out0 = v$COUT_998_out0;
assign v$RD_6030_out0 = v$CIN_9888_out0;
assign v$RD_6494_out0 = v$CIN_10112_out0;
assign v$G1_7885_out0 = ((v$RD_6030_out0 && !v$RM_11470_out0) || (!v$RD_6030_out0) && v$RM_11470_out0);
assign v$G1_8349_out0 = ((v$RD_6494_out0 && !v$RM_11934_out0) || (!v$RD_6494_out0) && v$RM_11934_out0);
assign v$G2_12421_out0 = v$RD_6030_out0 && v$RM_11470_out0;
assign v$G2_12885_out0 = v$RD_6494_out0 && v$RM_11934_out0;
assign v$CARRY_5030_out0 = v$G2_12421_out0;
assign v$CARRY_5494_out0 = v$G2_12885_out0;
assign v$S_9031_out0 = v$G1_7885_out0;
assign v$S_9495_out0 = v$G1_8349_out0;
assign v$S_1299_out0 = v$S_9031_out0;
assign v$S_1523_out0 = v$S_9495_out0;
assign v$G1_4075_out0 = v$CARRY_5030_out0 || v$CARRY_5029_out0;
assign v$G1_4299_out0 = v$CARRY_5494_out0 || v$CARRY_5493_out0;
assign v$COUT_767_out0 = v$G1_4075_out0;
assign v$COUT_991_out0 = v$G1_4299_out0;
assign v$_6931_out0 = { v$_4754_out0,v$S_1299_out0 };
assign v$_6946_out0 = { v$_4769_out0,v$S_1523_out0 };
assign v$CIN_9889_out0 = v$COUT_767_out0;
assign v$CIN_10113_out0 = v$COUT_991_out0;
assign v$RD_6032_out0 = v$CIN_9889_out0;
assign v$RD_6496_out0 = v$CIN_10113_out0;
assign v$G1_7887_out0 = ((v$RD_6032_out0 && !v$RM_11472_out0) || (!v$RD_6032_out0) && v$RM_11472_out0);
assign v$G1_8351_out0 = ((v$RD_6496_out0 && !v$RM_11936_out0) || (!v$RD_6496_out0) && v$RM_11936_out0);
assign v$G2_12423_out0 = v$RD_6032_out0 && v$RM_11472_out0;
assign v$G2_12887_out0 = v$RD_6496_out0 && v$RM_11936_out0;
assign v$CARRY_5032_out0 = v$G2_12423_out0;
assign v$CARRY_5496_out0 = v$G2_12887_out0;
assign v$S_9033_out0 = v$G1_7887_out0;
assign v$S_9497_out0 = v$G1_8351_out0;
assign v$S_1300_out0 = v$S_9033_out0;
assign v$S_1524_out0 = v$S_9497_out0;
assign v$G1_4076_out0 = v$CARRY_5032_out0 || v$CARRY_5031_out0;
assign v$G1_4300_out0 = v$CARRY_5496_out0 || v$CARRY_5495_out0;
assign v$COUT_768_out0 = v$G1_4076_out0;
assign v$COUT_992_out0 = v$G1_4300_out0;
assign v$_5807_out0 = { v$_6931_out0,v$S_1300_out0 };
assign v$_5822_out0 = { v$_6946_out0,v$S_1524_out0 };
assign v$CIN_9894_out0 = v$COUT_768_out0;
assign v$CIN_10118_out0 = v$COUT_992_out0;
assign v$RD_6042_out0 = v$CIN_9894_out0;
assign v$RD_6506_out0 = v$CIN_10118_out0;
assign v$G1_7897_out0 = ((v$RD_6042_out0 && !v$RM_11482_out0) || (!v$RD_6042_out0) && v$RM_11482_out0);
assign v$G1_8361_out0 = ((v$RD_6506_out0 && !v$RM_11946_out0) || (!v$RD_6506_out0) && v$RM_11946_out0);
assign v$G2_12433_out0 = v$RD_6042_out0 && v$RM_11482_out0;
assign v$G2_12897_out0 = v$RD_6506_out0 && v$RM_11946_out0;
assign v$CARRY_5042_out0 = v$G2_12433_out0;
assign v$CARRY_5506_out0 = v$G2_12897_out0;
assign v$S_9043_out0 = v$G1_7897_out0;
assign v$S_9507_out0 = v$G1_8361_out0;
assign v$S_1305_out0 = v$S_9043_out0;
assign v$S_1529_out0 = v$S_9507_out0;
assign v$G1_4081_out0 = v$CARRY_5042_out0 || v$CARRY_5041_out0;
assign v$G1_4305_out0 = v$CARRY_5506_out0 || v$CARRY_5505_out0;
assign v$COUT_773_out0 = v$G1_4081_out0;
assign v$COUT_997_out0 = v$G1_4305_out0;
assign v$_2031_out0 = { v$_5807_out0,v$S_1305_out0 };
assign v$_2046_out0 = { v$_5822_out0,v$S_1529_out0 };
assign v$CIN_9882_out0 = v$COUT_773_out0;
assign v$CIN_10106_out0 = v$COUT_997_out0;
assign v$RD_6017_out0 = v$CIN_9882_out0;
assign v$RD_6481_out0 = v$CIN_10106_out0;
assign v$G1_7872_out0 = ((v$RD_6017_out0 && !v$RM_11457_out0) || (!v$RD_6017_out0) && v$RM_11457_out0);
assign v$G1_8336_out0 = ((v$RD_6481_out0 && !v$RM_11921_out0) || (!v$RD_6481_out0) && v$RM_11921_out0);
assign v$G2_12408_out0 = v$RD_6017_out0 && v$RM_11457_out0;
assign v$G2_12872_out0 = v$RD_6481_out0 && v$RM_11921_out0;
assign v$CARRY_5017_out0 = v$G2_12408_out0;
assign v$CARRY_5481_out0 = v$G2_12872_out0;
assign v$S_9018_out0 = v$G1_7872_out0;
assign v$S_9482_out0 = v$G1_8336_out0;
assign v$S_1293_out0 = v$S_9018_out0;
assign v$S_1517_out0 = v$S_9482_out0;
assign v$G1_4069_out0 = v$CARRY_5017_out0 || v$CARRY_5016_out0;
assign v$G1_4293_out0 = v$CARRY_5481_out0 || v$CARRY_5480_out0;
assign v$COUT_761_out0 = v$G1_4069_out0;
assign v$COUT_985_out0 = v$G1_4293_out0;
assign v$_2798_out0 = { v$_2031_out0,v$S_1293_out0 };
assign v$_2813_out0 = { v$_2046_out0,v$S_1517_out0 };
assign v$CIN_9887_out0 = v$COUT_761_out0;
assign v$CIN_10111_out0 = v$COUT_985_out0;
assign v$RD_6027_out0 = v$CIN_9887_out0;
assign v$RD_6491_out0 = v$CIN_10111_out0;
assign v$G1_7882_out0 = ((v$RD_6027_out0 && !v$RM_11467_out0) || (!v$RD_6027_out0) && v$RM_11467_out0);
assign v$G1_8346_out0 = ((v$RD_6491_out0 && !v$RM_11931_out0) || (!v$RD_6491_out0) && v$RM_11931_out0);
assign v$G2_12418_out0 = v$RD_6027_out0 && v$RM_11467_out0;
assign v$G2_12882_out0 = v$RD_6491_out0 && v$RM_11931_out0;
assign v$CARRY_5027_out0 = v$G2_12418_out0;
assign v$CARRY_5491_out0 = v$G2_12882_out0;
assign v$S_9028_out0 = v$G1_7882_out0;
assign v$S_9492_out0 = v$G1_8346_out0;
assign v$S_1298_out0 = v$S_9028_out0;
assign v$S_1522_out0 = v$S_9492_out0;
assign v$G1_4074_out0 = v$CARRY_5027_out0 || v$CARRY_5026_out0;
assign v$G1_4298_out0 = v$CARRY_5491_out0 || v$CARRY_5490_out0;
assign v$COUT_766_out0 = v$G1_4074_out0;
assign v$COUT_990_out0 = v$G1_4298_out0;
assign v$_1830_out0 = { v$_2798_out0,v$S_1298_out0 };
assign v$_1845_out0 = { v$_2813_out0,v$S_1522_out0 };
assign v$CIN_9883_out0 = v$COUT_766_out0;
assign v$CIN_10107_out0 = v$COUT_990_out0;
assign v$RD_6019_out0 = v$CIN_9883_out0;
assign v$RD_6483_out0 = v$CIN_10107_out0;
assign v$G1_7874_out0 = ((v$RD_6019_out0 && !v$RM_11459_out0) || (!v$RD_6019_out0) && v$RM_11459_out0);
assign v$G1_8338_out0 = ((v$RD_6483_out0 && !v$RM_11923_out0) || (!v$RD_6483_out0) && v$RM_11923_out0);
assign v$G2_12410_out0 = v$RD_6019_out0 && v$RM_11459_out0;
assign v$G2_12874_out0 = v$RD_6483_out0 && v$RM_11923_out0;
assign v$CARRY_5019_out0 = v$G2_12410_out0;
assign v$CARRY_5483_out0 = v$G2_12874_out0;
assign v$S_9020_out0 = v$G1_7874_out0;
assign v$S_9484_out0 = v$G1_8338_out0;
assign v$S_1294_out0 = v$S_9020_out0;
assign v$S_1518_out0 = v$S_9484_out0;
assign v$G1_4070_out0 = v$CARRY_5019_out0 || v$CARRY_5018_out0;
assign v$G1_4294_out0 = v$CARRY_5483_out0 || v$CARRY_5482_out0;
assign v$COUT_762_out0 = v$G1_4070_out0;
assign v$COUT_986_out0 = v$G1_4294_out0;
assign v$_4554_out0 = { v$_1830_out0,v$S_1294_out0 };
assign v$_4569_out0 = { v$_1845_out0,v$S_1518_out0 };
assign v$RM_3431_out0 = v$COUT_762_out0;
assign v$RM_3655_out0 = v$COUT_986_out0;
assign v$RM_11460_out0 = v$RM_3431_out0;
assign v$RM_11924_out0 = v$RM_3655_out0;
assign v$G1_7875_out0 = ((v$RD_6020_out0 && !v$RM_11460_out0) || (!v$RD_6020_out0) && v$RM_11460_out0);
assign v$G1_8339_out0 = ((v$RD_6484_out0 && !v$RM_11924_out0) || (!v$RD_6484_out0) && v$RM_11924_out0);
assign v$G2_12411_out0 = v$RD_6020_out0 && v$RM_11460_out0;
assign v$G2_12875_out0 = v$RD_6484_out0 && v$RM_11924_out0;
assign v$CARRY_5020_out0 = v$G2_12411_out0;
assign v$CARRY_5484_out0 = v$G2_12875_out0;
assign v$S_9021_out0 = v$G1_7875_out0;
assign v$S_9485_out0 = v$G1_8339_out0;
assign v$RM_11461_out0 = v$S_9021_out0;
assign v$RM_11925_out0 = v$S_9485_out0;
assign v$G1_7876_out0 = ((v$RD_6021_out0 && !v$RM_11461_out0) || (!v$RD_6021_out0) && v$RM_11461_out0);
assign v$G1_8340_out0 = ((v$RD_6485_out0 && !v$RM_11925_out0) || (!v$RD_6485_out0) && v$RM_11925_out0);
assign v$G2_12412_out0 = v$RD_6021_out0 && v$RM_11461_out0;
assign v$G2_12876_out0 = v$RD_6485_out0 && v$RM_11925_out0;
assign v$CARRY_5021_out0 = v$G2_12412_out0;
assign v$CARRY_5485_out0 = v$G2_12876_out0;
assign v$S_9022_out0 = v$G1_7876_out0;
assign v$S_9486_out0 = v$G1_8340_out0;
assign v$S_1295_out0 = v$S_9022_out0;
assign v$S_1519_out0 = v$S_9486_out0;
assign v$G1_4071_out0 = v$CARRY_5021_out0 || v$CARRY_5020_out0;
assign v$G1_4295_out0 = v$CARRY_5485_out0 || v$CARRY_5484_out0;
assign v$COUT_763_out0 = v$G1_4071_out0;
assign v$COUT_987_out0 = v$G1_4295_out0;
assign v$_10656_out0 = { v$_4554_out0,v$S_1295_out0 };
assign v$_10671_out0 = { v$_4569_out0,v$S_1519_out0 };
assign v$_10951_out0 = { v$_10656_out0,v$COUT_763_out0 };
assign v$_10966_out0 = { v$_10671_out0,v$COUT_987_out0 };
assign v$COUT_10921_out0 = v$_10951_out0;
assign v$COUT_10936_out0 = v$_10966_out0;
assign v$CIN_2358_out0 = v$COUT_10921_out0;
assign v$CIN_2373_out0 = v$COUT_10936_out0;
assign v$_471_out0 = v$CIN_2358_out0[8:8];
assign v$_486_out0 = v$CIN_2373_out0[8:8];
assign v$_1776_out0 = v$CIN_2358_out0[6:6];
assign v$_1791_out0 = v$CIN_2373_out0[6:6];
assign v$_2158_out0 = v$CIN_2358_out0[3:3];
assign v$_2173_out0 = v$CIN_2373_out0[3:3];
assign v$_2197_out0 = v$CIN_2358_out0[15:15];
assign v$_2211_out0 = v$CIN_2373_out0[15:15];
assign v$_2505_out0 = v$CIN_2358_out0[0:0];
assign v$_2520_out0 = v$CIN_2373_out0[0:0];
assign v$_3054_out0 = v$CIN_2358_out0[9:9];
assign v$_3069_out0 = v$CIN_2373_out0[9:9];
assign v$_3088_out0 = v$CIN_2358_out0[2:2];
assign v$_3103_out0 = v$CIN_2373_out0[2:2];
assign v$_3142_out0 = v$CIN_2358_out0[7:7];
assign v$_3157_out0 = v$CIN_2373_out0[7:7];
assign v$_3826_out0 = v$CIN_2358_out0[1:1];
assign v$_3841_out0 = v$CIN_2373_out0[1:1];
assign v$_3864_out0 = v$CIN_2358_out0[10:10];
assign v$_3879_out0 = v$CIN_2373_out0[10:10];
assign v$_6803_out0 = v$CIN_2358_out0[11:11];
assign v$_6818_out0 = v$CIN_2373_out0[11:11];
assign v$_7647_out0 = v$CIN_2358_out0[12:12];
assign v$_7662_out0 = v$CIN_2373_out0[12:12];
assign v$_8702_out0 = v$CIN_2358_out0[13:13];
assign v$_8717_out0 = v$CIN_2373_out0[13:13];
assign v$_8772_out0 = v$CIN_2358_out0[14:14];
assign v$_8787_out0 = v$CIN_2373_out0[14:14];
assign v$_10722_out0 = v$CIN_2358_out0[5:5];
assign v$_10737_out0 = v$CIN_2373_out0[5:5];
assign v$_13451_out0 = v$CIN_2358_out0[4:4];
assign v$_13466_out0 = v$CIN_2373_out0[4:4];
assign v$RM_3399_out0 = v$_7647_out0;
assign v$RM_3400_out0 = v$_8772_out0;
assign v$RM_3402_out0 = v$_10722_out0;
assign v$RM_3403_out0 = v$_13451_out0;
assign v$RM_3404_out0 = v$_8702_out0;
assign v$RM_3405_out0 = v$_3054_out0;
assign v$RM_3406_out0 = v$_3864_out0;
assign v$RM_3407_out0 = v$_3826_out0;
assign v$RM_3408_out0 = v$_2158_out0;
assign v$RM_3409_out0 = v$_1776_out0;
assign v$RM_3410_out0 = v$_3142_out0;
assign v$RM_3411_out0 = v$_6803_out0;
assign v$RM_3412_out0 = v$_471_out0;
assign v$RM_3413_out0 = v$_3088_out0;
assign v$RM_3623_out0 = v$_7662_out0;
assign v$RM_3624_out0 = v$_8787_out0;
assign v$RM_3626_out0 = v$_10737_out0;
assign v$RM_3627_out0 = v$_13466_out0;
assign v$RM_3628_out0 = v$_8717_out0;
assign v$RM_3629_out0 = v$_3069_out0;
assign v$RM_3630_out0 = v$_3879_out0;
assign v$RM_3631_out0 = v$_3841_out0;
assign v$RM_3632_out0 = v$_2173_out0;
assign v$RM_3633_out0 = v$_1791_out0;
assign v$RM_3634_out0 = v$_3157_out0;
assign v$RM_3635_out0 = v$_6818_out0;
assign v$RM_3636_out0 = v$_486_out0;
assign v$RM_3637_out0 = v$_3103_out0;
assign v$CIN_9854_out0 = v$_2197_out0;
assign v$CIN_10078_out0 = v$_2211_out0;
assign v$RM_11406_out0 = v$_2505_out0;
assign v$RM_11870_out0 = v$_2520_out0;
assign v$RD_5959_out0 = v$CIN_9854_out0;
assign v$RD_6423_out0 = v$CIN_10078_out0;
assign v$G1_7821_out0 = ((v$RD_5966_out0 && !v$RM_11406_out0) || (!v$RD_5966_out0) && v$RM_11406_out0);
assign v$G1_8285_out0 = ((v$RD_6430_out0 && !v$RM_11870_out0) || (!v$RD_6430_out0) && v$RM_11870_out0);
assign v$RM_11394_out0 = v$RM_3399_out0;
assign v$RM_11396_out0 = v$RM_3400_out0;
assign v$RM_11400_out0 = v$RM_3402_out0;
assign v$RM_11402_out0 = v$RM_3403_out0;
assign v$RM_11404_out0 = v$RM_3404_out0;
assign v$RM_11407_out0 = v$RM_3405_out0;
assign v$RM_11409_out0 = v$RM_3406_out0;
assign v$RM_11411_out0 = v$RM_3407_out0;
assign v$RM_11413_out0 = v$RM_3408_out0;
assign v$RM_11415_out0 = v$RM_3409_out0;
assign v$RM_11417_out0 = v$RM_3410_out0;
assign v$RM_11419_out0 = v$RM_3411_out0;
assign v$RM_11421_out0 = v$RM_3412_out0;
assign v$RM_11423_out0 = v$RM_3413_out0;
assign v$RM_11858_out0 = v$RM_3623_out0;
assign v$RM_11860_out0 = v$RM_3624_out0;
assign v$RM_11864_out0 = v$RM_3626_out0;
assign v$RM_11866_out0 = v$RM_3627_out0;
assign v$RM_11868_out0 = v$RM_3628_out0;
assign v$RM_11871_out0 = v$RM_3629_out0;
assign v$RM_11873_out0 = v$RM_3630_out0;
assign v$RM_11875_out0 = v$RM_3631_out0;
assign v$RM_11877_out0 = v$RM_3632_out0;
assign v$RM_11879_out0 = v$RM_3633_out0;
assign v$RM_11881_out0 = v$RM_3634_out0;
assign v$RM_11883_out0 = v$RM_3635_out0;
assign v$RM_11885_out0 = v$RM_3636_out0;
assign v$RM_11887_out0 = v$RM_3637_out0;
assign v$G2_12357_out0 = v$RD_5966_out0 && v$RM_11406_out0;
assign v$G2_12821_out0 = v$RD_6430_out0 && v$RM_11870_out0;
assign v$CARRY_4966_out0 = v$G2_12357_out0;
assign v$CARRY_5430_out0 = v$G2_12821_out0;
assign v$G1_7809_out0 = ((v$RD_5954_out0 && !v$RM_11394_out0) || (!v$RD_5954_out0) && v$RM_11394_out0);
assign v$G1_7811_out0 = ((v$RD_5956_out0 && !v$RM_11396_out0) || (!v$RD_5956_out0) && v$RM_11396_out0);
assign v$G1_7815_out0 = ((v$RD_5960_out0 && !v$RM_11400_out0) || (!v$RD_5960_out0) && v$RM_11400_out0);
assign v$G1_7817_out0 = ((v$RD_5962_out0 && !v$RM_11402_out0) || (!v$RD_5962_out0) && v$RM_11402_out0);
assign v$G1_7819_out0 = ((v$RD_5964_out0 && !v$RM_11404_out0) || (!v$RD_5964_out0) && v$RM_11404_out0);
assign v$G1_7822_out0 = ((v$RD_5967_out0 && !v$RM_11407_out0) || (!v$RD_5967_out0) && v$RM_11407_out0);
assign v$G1_7824_out0 = ((v$RD_5969_out0 && !v$RM_11409_out0) || (!v$RD_5969_out0) && v$RM_11409_out0);
assign v$G1_7826_out0 = ((v$RD_5971_out0 && !v$RM_11411_out0) || (!v$RD_5971_out0) && v$RM_11411_out0);
assign v$G1_7828_out0 = ((v$RD_5973_out0 && !v$RM_11413_out0) || (!v$RD_5973_out0) && v$RM_11413_out0);
assign v$G1_7830_out0 = ((v$RD_5975_out0 && !v$RM_11415_out0) || (!v$RD_5975_out0) && v$RM_11415_out0);
assign v$G1_7832_out0 = ((v$RD_5977_out0 && !v$RM_11417_out0) || (!v$RD_5977_out0) && v$RM_11417_out0);
assign v$G1_7834_out0 = ((v$RD_5979_out0 && !v$RM_11419_out0) || (!v$RD_5979_out0) && v$RM_11419_out0);
assign v$G1_7836_out0 = ((v$RD_5981_out0 && !v$RM_11421_out0) || (!v$RD_5981_out0) && v$RM_11421_out0);
assign v$G1_7838_out0 = ((v$RD_5983_out0 && !v$RM_11423_out0) || (!v$RD_5983_out0) && v$RM_11423_out0);
assign v$G1_8273_out0 = ((v$RD_6418_out0 && !v$RM_11858_out0) || (!v$RD_6418_out0) && v$RM_11858_out0);
assign v$G1_8275_out0 = ((v$RD_6420_out0 && !v$RM_11860_out0) || (!v$RD_6420_out0) && v$RM_11860_out0);
assign v$G1_8279_out0 = ((v$RD_6424_out0 && !v$RM_11864_out0) || (!v$RD_6424_out0) && v$RM_11864_out0);
assign v$G1_8281_out0 = ((v$RD_6426_out0 && !v$RM_11866_out0) || (!v$RD_6426_out0) && v$RM_11866_out0);
assign v$G1_8283_out0 = ((v$RD_6428_out0 && !v$RM_11868_out0) || (!v$RD_6428_out0) && v$RM_11868_out0);
assign v$G1_8286_out0 = ((v$RD_6431_out0 && !v$RM_11871_out0) || (!v$RD_6431_out0) && v$RM_11871_out0);
assign v$G1_8288_out0 = ((v$RD_6433_out0 && !v$RM_11873_out0) || (!v$RD_6433_out0) && v$RM_11873_out0);
assign v$G1_8290_out0 = ((v$RD_6435_out0 && !v$RM_11875_out0) || (!v$RD_6435_out0) && v$RM_11875_out0);
assign v$G1_8292_out0 = ((v$RD_6437_out0 && !v$RM_11877_out0) || (!v$RD_6437_out0) && v$RM_11877_out0);
assign v$G1_8294_out0 = ((v$RD_6439_out0 && !v$RM_11879_out0) || (!v$RD_6439_out0) && v$RM_11879_out0);
assign v$G1_8296_out0 = ((v$RD_6441_out0 && !v$RM_11881_out0) || (!v$RD_6441_out0) && v$RM_11881_out0);
assign v$G1_8298_out0 = ((v$RD_6443_out0 && !v$RM_11883_out0) || (!v$RD_6443_out0) && v$RM_11883_out0);
assign v$G1_8300_out0 = ((v$RD_6445_out0 && !v$RM_11885_out0) || (!v$RD_6445_out0) && v$RM_11885_out0);
assign v$G1_8302_out0 = ((v$RD_6447_out0 && !v$RM_11887_out0) || (!v$RD_6447_out0) && v$RM_11887_out0);
assign v$S_8967_out0 = v$G1_7821_out0;
assign v$S_9431_out0 = v$G1_8285_out0;
assign v$G2_12345_out0 = v$RD_5954_out0 && v$RM_11394_out0;
assign v$G2_12347_out0 = v$RD_5956_out0 && v$RM_11396_out0;
assign v$G2_12351_out0 = v$RD_5960_out0 && v$RM_11400_out0;
assign v$G2_12353_out0 = v$RD_5962_out0 && v$RM_11402_out0;
assign v$G2_12355_out0 = v$RD_5964_out0 && v$RM_11404_out0;
assign v$G2_12358_out0 = v$RD_5967_out0 && v$RM_11407_out0;
assign v$G2_12360_out0 = v$RD_5969_out0 && v$RM_11409_out0;
assign v$G2_12362_out0 = v$RD_5971_out0 && v$RM_11411_out0;
assign v$G2_12364_out0 = v$RD_5973_out0 && v$RM_11413_out0;
assign v$G2_12366_out0 = v$RD_5975_out0 && v$RM_11415_out0;
assign v$G2_12368_out0 = v$RD_5977_out0 && v$RM_11417_out0;
assign v$G2_12370_out0 = v$RD_5979_out0 && v$RM_11419_out0;
assign v$G2_12372_out0 = v$RD_5981_out0 && v$RM_11421_out0;
assign v$G2_12374_out0 = v$RD_5983_out0 && v$RM_11423_out0;
assign v$G2_12809_out0 = v$RD_6418_out0 && v$RM_11858_out0;
assign v$G2_12811_out0 = v$RD_6420_out0 && v$RM_11860_out0;
assign v$G2_12815_out0 = v$RD_6424_out0 && v$RM_11864_out0;
assign v$G2_12817_out0 = v$RD_6426_out0 && v$RM_11866_out0;
assign v$G2_12819_out0 = v$RD_6428_out0 && v$RM_11868_out0;
assign v$G2_12822_out0 = v$RD_6431_out0 && v$RM_11871_out0;
assign v$G2_12824_out0 = v$RD_6433_out0 && v$RM_11873_out0;
assign v$G2_12826_out0 = v$RD_6435_out0 && v$RM_11875_out0;
assign v$G2_12828_out0 = v$RD_6437_out0 && v$RM_11877_out0;
assign v$G2_12830_out0 = v$RD_6439_out0 && v$RM_11879_out0;
assign v$G2_12832_out0 = v$RD_6441_out0 && v$RM_11881_out0;
assign v$G2_12834_out0 = v$RD_6443_out0 && v$RM_11883_out0;
assign v$G2_12836_out0 = v$RD_6445_out0 && v$RM_11885_out0;
assign v$G2_12838_out0 = v$RD_6447_out0 && v$RM_11887_out0;
assign v$S_4668_out0 = v$S_8967_out0;
assign v$S_4683_out0 = v$S_9431_out0;
assign v$CARRY_4954_out0 = v$G2_12345_out0;
assign v$CARRY_4956_out0 = v$G2_12347_out0;
assign v$CARRY_4960_out0 = v$G2_12351_out0;
assign v$CARRY_4962_out0 = v$G2_12353_out0;
assign v$CARRY_4964_out0 = v$G2_12355_out0;
assign v$CARRY_4967_out0 = v$G2_12358_out0;
assign v$CARRY_4969_out0 = v$G2_12360_out0;
assign v$CARRY_4971_out0 = v$G2_12362_out0;
assign v$CARRY_4973_out0 = v$G2_12364_out0;
assign v$CARRY_4975_out0 = v$G2_12366_out0;
assign v$CARRY_4977_out0 = v$G2_12368_out0;
assign v$CARRY_4979_out0 = v$G2_12370_out0;
assign v$CARRY_4981_out0 = v$G2_12372_out0;
assign v$CARRY_4983_out0 = v$G2_12374_out0;
assign v$CARRY_5418_out0 = v$G2_12809_out0;
assign v$CARRY_5420_out0 = v$G2_12811_out0;
assign v$CARRY_5424_out0 = v$G2_12815_out0;
assign v$CARRY_5426_out0 = v$G2_12817_out0;
assign v$CARRY_5428_out0 = v$G2_12819_out0;
assign v$CARRY_5431_out0 = v$G2_12822_out0;
assign v$CARRY_5433_out0 = v$G2_12824_out0;
assign v$CARRY_5435_out0 = v$G2_12826_out0;
assign v$CARRY_5437_out0 = v$G2_12828_out0;
assign v$CARRY_5439_out0 = v$G2_12830_out0;
assign v$CARRY_5441_out0 = v$G2_12832_out0;
assign v$CARRY_5443_out0 = v$G2_12834_out0;
assign v$CARRY_5445_out0 = v$G2_12836_out0;
assign v$CARRY_5447_out0 = v$G2_12838_out0;
assign v$S_8955_out0 = v$G1_7809_out0;
assign v$S_8957_out0 = v$G1_7811_out0;
assign v$S_8961_out0 = v$G1_7815_out0;
assign v$S_8963_out0 = v$G1_7817_out0;
assign v$S_8965_out0 = v$G1_7819_out0;
assign v$S_8968_out0 = v$G1_7822_out0;
assign v$S_8970_out0 = v$G1_7824_out0;
assign v$S_8972_out0 = v$G1_7826_out0;
assign v$S_8974_out0 = v$G1_7828_out0;
assign v$S_8976_out0 = v$G1_7830_out0;
assign v$S_8978_out0 = v$G1_7832_out0;
assign v$S_8980_out0 = v$G1_7834_out0;
assign v$S_8982_out0 = v$G1_7836_out0;
assign v$S_8984_out0 = v$G1_7838_out0;
assign v$S_9419_out0 = v$G1_8273_out0;
assign v$S_9421_out0 = v$G1_8275_out0;
assign v$S_9425_out0 = v$G1_8279_out0;
assign v$S_9427_out0 = v$G1_8281_out0;
assign v$S_9429_out0 = v$G1_8283_out0;
assign v$S_9432_out0 = v$G1_8286_out0;
assign v$S_9434_out0 = v$G1_8288_out0;
assign v$S_9436_out0 = v$G1_8290_out0;
assign v$S_9438_out0 = v$G1_8292_out0;
assign v$S_9440_out0 = v$G1_8294_out0;
assign v$S_9442_out0 = v$G1_8296_out0;
assign v$S_9444_out0 = v$G1_8298_out0;
assign v$S_9446_out0 = v$G1_8300_out0;
assign v$S_9448_out0 = v$G1_8302_out0;
assign v$CIN_9860_out0 = v$CARRY_4966_out0;
assign v$CIN_10084_out0 = v$CARRY_5430_out0;
assign v$_2439_out0 = { v$_2191_out0,v$S_4668_out0 };
assign v$_2440_out0 = { v$_2192_out0,v$S_4683_out0 };
assign v$RD_5972_out0 = v$CIN_9860_out0;
assign v$RD_6436_out0 = v$CIN_10084_out0;
assign v$RM_11395_out0 = v$S_8955_out0;
assign v$RM_11397_out0 = v$S_8957_out0;
assign v$RM_11401_out0 = v$S_8961_out0;
assign v$RM_11403_out0 = v$S_8963_out0;
assign v$RM_11405_out0 = v$S_8965_out0;
assign v$RM_11408_out0 = v$S_8968_out0;
assign v$RM_11410_out0 = v$S_8970_out0;
assign v$RM_11412_out0 = v$S_8972_out0;
assign v$RM_11414_out0 = v$S_8974_out0;
assign v$RM_11416_out0 = v$S_8976_out0;
assign v$RM_11418_out0 = v$S_8978_out0;
assign v$RM_11420_out0 = v$S_8980_out0;
assign v$RM_11422_out0 = v$S_8982_out0;
assign v$RM_11424_out0 = v$S_8984_out0;
assign v$RM_11859_out0 = v$S_9419_out0;
assign v$RM_11861_out0 = v$S_9421_out0;
assign v$RM_11865_out0 = v$S_9425_out0;
assign v$RM_11867_out0 = v$S_9427_out0;
assign v$RM_11869_out0 = v$S_9429_out0;
assign v$RM_11872_out0 = v$S_9432_out0;
assign v$RM_11874_out0 = v$S_9434_out0;
assign v$RM_11876_out0 = v$S_9436_out0;
assign v$RM_11878_out0 = v$S_9438_out0;
assign v$RM_11880_out0 = v$S_9440_out0;
assign v$RM_11882_out0 = v$S_9442_out0;
assign v$RM_11884_out0 = v$S_9444_out0;
assign v$RM_11886_out0 = v$S_9446_out0;
assign v$RM_11888_out0 = v$S_9448_out0;
assign v$G1_7827_out0 = ((v$RD_5972_out0 && !v$RM_11412_out0) || (!v$RD_5972_out0) && v$RM_11412_out0);
assign v$G1_8291_out0 = ((v$RD_6436_out0 && !v$RM_11876_out0) || (!v$RD_6436_out0) && v$RM_11876_out0);
assign v$G2_12363_out0 = v$RD_5972_out0 && v$RM_11412_out0;
assign v$G2_12827_out0 = v$RD_6436_out0 && v$RM_11876_out0;
assign v$CARRY_4972_out0 = v$G2_12363_out0;
assign v$CARRY_5436_out0 = v$G2_12827_out0;
assign v$S_8973_out0 = v$G1_7827_out0;
assign v$S_9437_out0 = v$G1_8291_out0;
assign v$S_1271_out0 = v$S_8973_out0;
assign v$S_1495_out0 = v$S_9437_out0;
assign v$G1_4047_out0 = v$CARRY_4972_out0 || v$CARRY_4971_out0;
assign v$G1_4271_out0 = v$CARRY_5436_out0 || v$CARRY_5435_out0;
assign v$COUT_739_out0 = v$G1_4047_out0;
assign v$COUT_963_out0 = v$G1_4271_out0;
assign v$CIN_9866_out0 = v$COUT_739_out0;
assign v$CIN_10090_out0 = v$COUT_963_out0;
assign v$RD_5984_out0 = v$CIN_9866_out0;
assign v$RD_6448_out0 = v$CIN_10090_out0;
assign v$G1_7839_out0 = ((v$RD_5984_out0 && !v$RM_11424_out0) || (!v$RD_5984_out0) && v$RM_11424_out0);
assign v$G1_8303_out0 = ((v$RD_6448_out0 && !v$RM_11888_out0) || (!v$RD_6448_out0) && v$RM_11888_out0);
assign v$G2_12375_out0 = v$RD_5984_out0 && v$RM_11424_out0;
assign v$G2_12839_out0 = v$RD_6448_out0 && v$RM_11888_out0;
assign v$CARRY_4984_out0 = v$G2_12375_out0;
assign v$CARRY_5448_out0 = v$G2_12839_out0;
assign v$S_8985_out0 = v$G1_7839_out0;
assign v$S_9449_out0 = v$G1_8303_out0;
assign v$S_1277_out0 = v$S_8985_out0;
assign v$S_1501_out0 = v$S_9449_out0;
assign v$G1_4053_out0 = v$CARRY_4984_out0 || v$CARRY_4983_out0;
assign v$G1_4277_out0 = v$CARRY_5448_out0 || v$CARRY_5447_out0;
assign v$COUT_745_out0 = v$G1_4053_out0;
assign v$COUT_969_out0 = v$G1_4277_out0;
assign v$_4785_out0 = { v$S_1271_out0,v$S_1277_out0 };
assign v$_4800_out0 = { v$S_1495_out0,v$S_1501_out0 };
assign v$CIN_9861_out0 = v$COUT_745_out0;
assign v$CIN_10085_out0 = v$COUT_969_out0;
assign v$RD_5974_out0 = v$CIN_9861_out0;
assign v$RD_6438_out0 = v$CIN_10085_out0;
assign v$G1_7829_out0 = ((v$RD_5974_out0 && !v$RM_11414_out0) || (!v$RD_5974_out0) && v$RM_11414_out0);
assign v$G1_8293_out0 = ((v$RD_6438_out0 && !v$RM_11878_out0) || (!v$RD_6438_out0) && v$RM_11878_out0);
assign v$G2_12365_out0 = v$RD_5974_out0 && v$RM_11414_out0;
assign v$G2_12829_out0 = v$RD_6438_out0 && v$RM_11878_out0;
assign v$CARRY_4974_out0 = v$G2_12365_out0;
assign v$CARRY_5438_out0 = v$G2_12829_out0;
assign v$S_8975_out0 = v$G1_7829_out0;
assign v$S_9439_out0 = v$G1_8293_out0;
assign v$S_1272_out0 = v$S_8975_out0;
assign v$S_1496_out0 = v$S_9439_out0;
assign v$G1_4048_out0 = v$CARRY_4974_out0 || v$CARRY_4973_out0;
assign v$G1_4272_out0 = v$CARRY_5438_out0 || v$CARRY_5437_out0;
assign v$COUT_740_out0 = v$G1_4048_out0;
assign v$COUT_964_out0 = v$G1_4272_out0;
assign v$_2555_out0 = { v$_4785_out0,v$S_1272_out0 };
assign v$_2570_out0 = { v$_4800_out0,v$S_1496_out0 };
assign v$CIN_9856_out0 = v$COUT_740_out0;
assign v$CIN_10080_out0 = v$COUT_964_out0;
assign v$RD_5963_out0 = v$CIN_9856_out0;
assign v$RD_6427_out0 = v$CIN_10080_out0;
assign v$G1_7818_out0 = ((v$RD_5963_out0 && !v$RM_11403_out0) || (!v$RD_5963_out0) && v$RM_11403_out0);
assign v$G1_8282_out0 = ((v$RD_6427_out0 && !v$RM_11867_out0) || (!v$RD_6427_out0) && v$RM_11867_out0);
assign v$G2_12354_out0 = v$RD_5963_out0 && v$RM_11403_out0;
assign v$G2_12818_out0 = v$RD_6427_out0 && v$RM_11867_out0;
assign v$CARRY_4963_out0 = v$G2_12354_out0;
assign v$CARRY_5427_out0 = v$G2_12818_out0;
assign v$S_8964_out0 = v$G1_7818_out0;
assign v$S_9428_out0 = v$G1_8282_out0;
assign v$S_1267_out0 = v$S_8964_out0;
assign v$S_1491_out0 = v$S_9428_out0;
assign v$G1_4043_out0 = v$CARRY_4963_out0 || v$CARRY_4962_out0;
assign v$G1_4267_out0 = v$CARRY_5427_out0 || v$CARRY_5426_out0;
assign v$COUT_735_out0 = v$G1_4043_out0;
assign v$COUT_959_out0 = v$G1_4267_out0;
assign v$_7035_out0 = { v$_2555_out0,v$S_1267_out0 };
assign v$_7050_out0 = { v$_2570_out0,v$S_1491_out0 };
assign v$CIN_9855_out0 = v$COUT_735_out0;
assign v$CIN_10079_out0 = v$COUT_959_out0;
assign v$RD_5961_out0 = v$CIN_9855_out0;
assign v$RD_6425_out0 = v$CIN_10079_out0;
assign v$G1_7816_out0 = ((v$RD_5961_out0 && !v$RM_11401_out0) || (!v$RD_5961_out0) && v$RM_11401_out0);
assign v$G1_8280_out0 = ((v$RD_6425_out0 && !v$RM_11865_out0) || (!v$RD_6425_out0) && v$RM_11865_out0);
assign v$G2_12352_out0 = v$RD_5961_out0 && v$RM_11401_out0;
assign v$G2_12816_out0 = v$RD_6425_out0 && v$RM_11865_out0;
assign v$CARRY_4961_out0 = v$G2_12352_out0;
assign v$CARRY_5425_out0 = v$G2_12816_out0;
assign v$S_8962_out0 = v$G1_7816_out0;
assign v$S_9426_out0 = v$G1_8280_out0;
assign v$S_1266_out0 = v$S_8962_out0;
assign v$S_1490_out0 = v$S_9426_out0;
assign v$G1_4042_out0 = v$CARRY_4961_out0 || v$CARRY_4960_out0;
assign v$G1_4266_out0 = v$CARRY_5425_out0 || v$CARRY_5424_out0;
assign v$COUT_734_out0 = v$G1_4042_out0;
assign v$COUT_958_out0 = v$G1_4266_out0;
assign v$_13521_out0 = { v$_7035_out0,v$S_1266_out0 };
assign v$_13536_out0 = { v$_7050_out0,v$S_1490_out0 };
assign v$CIN_9862_out0 = v$COUT_734_out0;
assign v$CIN_10086_out0 = v$COUT_958_out0;
assign v$RD_5976_out0 = v$CIN_9862_out0;
assign v$RD_6440_out0 = v$CIN_10086_out0;
assign v$G1_7831_out0 = ((v$RD_5976_out0 && !v$RM_11416_out0) || (!v$RD_5976_out0) && v$RM_11416_out0);
assign v$G1_8295_out0 = ((v$RD_6440_out0 && !v$RM_11880_out0) || (!v$RD_6440_out0) && v$RM_11880_out0);
assign v$G2_12367_out0 = v$RD_5976_out0 && v$RM_11416_out0;
assign v$G2_12831_out0 = v$RD_6440_out0 && v$RM_11880_out0;
assign v$CARRY_4976_out0 = v$G2_12367_out0;
assign v$CARRY_5440_out0 = v$G2_12831_out0;
assign v$S_8977_out0 = v$G1_7831_out0;
assign v$S_9441_out0 = v$G1_8295_out0;
assign v$S_1273_out0 = v$S_8977_out0;
assign v$S_1497_out0 = v$S_9441_out0;
assign v$G1_4049_out0 = v$CARRY_4976_out0 || v$CARRY_4975_out0;
assign v$G1_4273_out0 = v$CARRY_5440_out0 || v$CARRY_5439_out0;
assign v$COUT_741_out0 = v$G1_4049_out0;
assign v$COUT_965_out0 = v$G1_4273_out0;
assign v$_3314_out0 = { v$_13521_out0,v$S_1273_out0 };
assign v$_3329_out0 = { v$_13536_out0,v$S_1497_out0 };
assign v$CIN_9863_out0 = v$COUT_741_out0;
assign v$CIN_10087_out0 = v$COUT_965_out0;
assign v$RD_5978_out0 = v$CIN_9863_out0;
assign v$RD_6442_out0 = v$CIN_10087_out0;
assign v$G1_7833_out0 = ((v$RD_5978_out0 && !v$RM_11418_out0) || (!v$RD_5978_out0) && v$RM_11418_out0);
assign v$G1_8297_out0 = ((v$RD_6442_out0 && !v$RM_11882_out0) || (!v$RD_6442_out0) && v$RM_11882_out0);
assign v$G2_12369_out0 = v$RD_5978_out0 && v$RM_11418_out0;
assign v$G2_12833_out0 = v$RD_6442_out0 && v$RM_11882_out0;
assign v$CARRY_4978_out0 = v$G2_12369_out0;
assign v$CARRY_5442_out0 = v$G2_12833_out0;
assign v$S_8979_out0 = v$G1_7833_out0;
assign v$S_9443_out0 = v$G1_8297_out0;
assign v$S_1274_out0 = v$S_8979_out0;
assign v$S_1498_out0 = v$S_9443_out0;
assign v$G1_4050_out0 = v$CARRY_4978_out0 || v$CARRY_4977_out0;
assign v$G1_4274_out0 = v$CARRY_5442_out0 || v$CARRY_5441_out0;
assign v$COUT_742_out0 = v$G1_4050_out0;
assign v$COUT_966_out0 = v$G1_4274_out0;
assign v$_7150_out0 = { v$_3314_out0,v$S_1274_out0 };
assign v$_7165_out0 = { v$_3329_out0,v$S_1498_out0 };
assign v$CIN_9865_out0 = v$COUT_742_out0;
assign v$CIN_10089_out0 = v$COUT_966_out0;
assign v$RD_5982_out0 = v$CIN_9865_out0;
assign v$RD_6446_out0 = v$CIN_10089_out0;
assign v$G1_7837_out0 = ((v$RD_5982_out0 && !v$RM_11422_out0) || (!v$RD_5982_out0) && v$RM_11422_out0);
assign v$G1_8301_out0 = ((v$RD_6446_out0 && !v$RM_11886_out0) || (!v$RD_6446_out0) && v$RM_11886_out0);
assign v$G2_12373_out0 = v$RD_5982_out0 && v$RM_11422_out0;
assign v$G2_12837_out0 = v$RD_6446_out0 && v$RM_11886_out0;
assign v$CARRY_4982_out0 = v$G2_12373_out0;
assign v$CARRY_5446_out0 = v$G2_12837_out0;
assign v$S_8983_out0 = v$G1_7837_out0;
assign v$S_9447_out0 = v$G1_8301_out0;
assign v$S_1276_out0 = v$S_8983_out0;
assign v$S_1500_out0 = v$S_9447_out0;
assign v$G1_4052_out0 = v$CARRY_4982_out0 || v$CARRY_4981_out0;
assign v$G1_4276_out0 = v$CARRY_5446_out0 || v$CARRY_5445_out0;
assign v$COUT_744_out0 = v$G1_4052_out0;
assign v$COUT_968_out0 = v$G1_4276_out0;
assign v$_4752_out0 = { v$_7150_out0,v$S_1276_out0 };
assign v$_4767_out0 = { v$_7165_out0,v$S_1500_out0 };
assign v$CIN_9858_out0 = v$COUT_744_out0;
assign v$CIN_10082_out0 = v$COUT_968_out0;
assign v$RD_5968_out0 = v$CIN_9858_out0;
assign v$RD_6432_out0 = v$CIN_10082_out0;
assign v$G1_7823_out0 = ((v$RD_5968_out0 && !v$RM_11408_out0) || (!v$RD_5968_out0) && v$RM_11408_out0);
assign v$G1_8287_out0 = ((v$RD_6432_out0 && !v$RM_11872_out0) || (!v$RD_6432_out0) && v$RM_11872_out0);
assign v$G2_12359_out0 = v$RD_5968_out0 && v$RM_11408_out0;
assign v$G2_12823_out0 = v$RD_6432_out0 && v$RM_11872_out0;
assign v$CARRY_4968_out0 = v$G2_12359_out0;
assign v$CARRY_5432_out0 = v$G2_12823_out0;
assign v$S_8969_out0 = v$G1_7823_out0;
assign v$S_9433_out0 = v$G1_8287_out0;
assign v$S_1269_out0 = v$S_8969_out0;
assign v$S_1493_out0 = v$S_9433_out0;
assign v$G1_4045_out0 = v$CARRY_4968_out0 || v$CARRY_4967_out0;
assign v$G1_4269_out0 = v$CARRY_5432_out0 || v$CARRY_5431_out0;
assign v$COUT_737_out0 = v$G1_4045_out0;
assign v$COUT_961_out0 = v$G1_4269_out0;
assign v$_6929_out0 = { v$_4752_out0,v$S_1269_out0 };
assign v$_6944_out0 = { v$_4767_out0,v$S_1493_out0 };
assign v$CIN_9859_out0 = v$COUT_737_out0;
assign v$CIN_10083_out0 = v$COUT_961_out0;
assign v$RD_5970_out0 = v$CIN_9859_out0;
assign v$RD_6434_out0 = v$CIN_10083_out0;
assign v$G1_7825_out0 = ((v$RD_5970_out0 && !v$RM_11410_out0) || (!v$RD_5970_out0) && v$RM_11410_out0);
assign v$G1_8289_out0 = ((v$RD_6434_out0 && !v$RM_11874_out0) || (!v$RD_6434_out0) && v$RM_11874_out0);
assign v$G2_12361_out0 = v$RD_5970_out0 && v$RM_11410_out0;
assign v$G2_12825_out0 = v$RD_6434_out0 && v$RM_11874_out0;
assign v$CARRY_4970_out0 = v$G2_12361_out0;
assign v$CARRY_5434_out0 = v$G2_12825_out0;
assign v$S_8971_out0 = v$G1_7825_out0;
assign v$S_9435_out0 = v$G1_8289_out0;
assign v$S_1270_out0 = v$S_8971_out0;
assign v$S_1494_out0 = v$S_9435_out0;
assign v$G1_4046_out0 = v$CARRY_4970_out0 || v$CARRY_4969_out0;
assign v$G1_4270_out0 = v$CARRY_5434_out0 || v$CARRY_5433_out0;
assign v$COUT_738_out0 = v$G1_4046_out0;
assign v$COUT_962_out0 = v$G1_4270_out0;
assign v$_5805_out0 = { v$_6929_out0,v$S_1270_out0 };
assign v$_5820_out0 = { v$_6944_out0,v$S_1494_out0 };
assign v$CIN_9864_out0 = v$COUT_738_out0;
assign v$CIN_10088_out0 = v$COUT_962_out0;
assign v$RD_5980_out0 = v$CIN_9864_out0;
assign v$RD_6444_out0 = v$CIN_10088_out0;
assign v$G1_7835_out0 = ((v$RD_5980_out0 && !v$RM_11420_out0) || (!v$RD_5980_out0) && v$RM_11420_out0);
assign v$G1_8299_out0 = ((v$RD_6444_out0 && !v$RM_11884_out0) || (!v$RD_6444_out0) && v$RM_11884_out0);
assign v$G2_12371_out0 = v$RD_5980_out0 && v$RM_11420_out0;
assign v$G2_12835_out0 = v$RD_6444_out0 && v$RM_11884_out0;
assign v$CARRY_4980_out0 = v$G2_12371_out0;
assign v$CARRY_5444_out0 = v$G2_12835_out0;
assign v$S_8981_out0 = v$G1_7835_out0;
assign v$S_9445_out0 = v$G1_8299_out0;
assign v$S_1275_out0 = v$S_8981_out0;
assign v$S_1499_out0 = v$S_9445_out0;
assign v$G1_4051_out0 = v$CARRY_4980_out0 || v$CARRY_4979_out0;
assign v$G1_4275_out0 = v$CARRY_5444_out0 || v$CARRY_5443_out0;
assign v$COUT_743_out0 = v$G1_4051_out0;
assign v$COUT_967_out0 = v$G1_4275_out0;
assign v$_2029_out0 = { v$_5805_out0,v$S_1275_out0 };
assign v$_2044_out0 = { v$_5820_out0,v$S_1499_out0 };
assign v$CIN_9852_out0 = v$COUT_743_out0;
assign v$CIN_10076_out0 = v$COUT_967_out0;
assign v$RD_5955_out0 = v$CIN_9852_out0;
assign v$RD_6419_out0 = v$CIN_10076_out0;
assign v$G1_7810_out0 = ((v$RD_5955_out0 && !v$RM_11395_out0) || (!v$RD_5955_out0) && v$RM_11395_out0);
assign v$G1_8274_out0 = ((v$RD_6419_out0 && !v$RM_11859_out0) || (!v$RD_6419_out0) && v$RM_11859_out0);
assign v$G2_12346_out0 = v$RD_5955_out0 && v$RM_11395_out0;
assign v$G2_12810_out0 = v$RD_6419_out0 && v$RM_11859_out0;
assign v$CARRY_4955_out0 = v$G2_12346_out0;
assign v$CARRY_5419_out0 = v$G2_12810_out0;
assign v$S_8956_out0 = v$G1_7810_out0;
assign v$S_9420_out0 = v$G1_8274_out0;
assign v$S_1263_out0 = v$S_8956_out0;
assign v$S_1487_out0 = v$S_9420_out0;
assign v$G1_4039_out0 = v$CARRY_4955_out0 || v$CARRY_4954_out0;
assign v$G1_4263_out0 = v$CARRY_5419_out0 || v$CARRY_5418_out0;
assign v$COUT_731_out0 = v$G1_4039_out0;
assign v$COUT_955_out0 = v$G1_4263_out0;
assign v$_2796_out0 = { v$_2029_out0,v$S_1263_out0 };
assign v$_2811_out0 = { v$_2044_out0,v$S_1487_out0 };
assign v$CIN_9857_out0 = v$COUT_731_out0;
assign v$CIN_10081_out0 = v$COUT_955_out0;
assign v$RD_5965_out0 = v$CIN_9857_out0;
assign v$RD_6429_out0 = v$CIN_10081_out0;
assign v$G1_7820_out0 = ((v$RD_5965_out0 && !v$RM_11405_out0) || (!v$RD_5965_out0) && v$RM_11405_out0);
assign v$G1_8284_out0 = ((v$RD_6429_out0 && !v$RM_11869_out0) || (!v$RD_6429_out0) && v$RM_11869_out0);
assign v$G2_12356_out0 = v$RD_5965_out0 && v$RM_11405_out0;
assign v$G2_12820_out0 = v$RD_6429_out0 && v$RM_11869_out0;
assign v$CARRY_4965_out0 = v$G2_12356_out0;
assign v$CARRY_5429_out0 = v$G2_12820_out0;
assign v$S_8966_out0 = v$G1_7820_out0;
assign v$S_9430_out0 = v$G1_8284_out0;
assign v$S_1268_out0 = v$S_8966_out0;
assign v$S_1492_out0 = v$S_9430_out0;
assign v$G1_4044_out0 = v$CARRY_4965_out0 || v$CARRY_4964_out0;
assign v$G1_4268_out0 = v$CARRY_5429_out0 || v$CARRY_5428_out0;
assign v$COUT_736_out0 = v$G1_4044_out0;
assign v$COUT_960_out0 = v$G1_4268_out0;
assign v$_1828_out0 = { v$_2796_out0,v$S_1268_out0 };
assign v$_1843_out0 = { v$_2811_out0,v$S_1492_out0 };
assign v$CIN_9853_out0 = v$COUT_736_out0;
assign v$CIN_10077_out0 = v$COUT_960_out0;
assign v$RD_5957_out0 = v$CIN_9853_out0;
assign v$RD_6421_out0 = v$CIN_10077_out0;
assign v$G1_7812_out0 = ((v$RD_5957_out0 && !v$RM_11397_out0) || (!v$RD_5957_out0) && v$RM_11397_out0);
assign v$G1_8276_out0 = ((v$RD_6421_out0 && !v$RM_11861_out0) || (!v$RD_6421_out0) && v$RM_11861_out0);
assign v$G2_12348_out0 = v$RD_5957_out0 && v$RM_11397_out0;
assign v$G2_12812_out0 = v$RD_6421_out0 && v$RM_11861_out0;
assign v$CARRY_4957_out0 = v$G2_12348_out0;
assign v$CARRY_5421_out0 = v$G2_12812_out0;
assign v$S_8958_out0 = v$G1_7812_out0;
assign v$S_9422_out0 = v$G1_8276_out0;
assign v$S_1264_out0 = v$S_8958_out0;
assign v$S_1488_out0 = v$S_9422_out0;
assign v$G1_4040_out0 = v$CARRY_4957_out0 || v$CARRY_4956_out0;
assign v$G1_4264_out0 = v$CARRY_5421_out0 || v$CARRY_5420_out0;
assign v$COUT_732_out0 = v$G1_4040_out0;
assign v$COUT_956_out0 = v$G1_4264_out0;
assign v$_4552_out0 = { v$_1828_out0,v$S_1264_out0 };
assign v$_4567_out0 = { v$_1843_out0,v$S_1488_out0 };
assign v$RM_3401_out0 = v$COUT_732_out0;
assign v$RM_3625_out0 = v$COUT_956_out0;
assign v$RM_11398_out0 = v$RM_3401_out0;
assign v$RM_11862_out0 = v$RM_3625_out0;
assign v$G1_7813_out0 = ((v$RD_5958_out0 && !v$RM_11398_out0) || (!v$RD_5958_out0) && v$RM_11398_out0);
assign v$G1_8277_out0 = ((v$RD_6422_out0 && !v$RM_11862_out0) || (!v$RD_6422_out0) && v$RM_11862_out0);
assign v$G2_12349_out0 = v$RD_5958_out0 && v$RM_11398_out0;
assign v$G2_12813_out0 = v$RD_6422_out0 && v$RM_11862_out0;
assign v$CARRY_4958_out0 = v$G2_12349_out0;
assign v$CARRY_5422_out0 = v$G2_12813_out0;
assign v$S_8959_out0 = v$G1_7813_out0;
assign v$S_9423_out0 = v$G1_8277_out0;
assign v$RM_11399_out0 = v$S_8959_out0;
assign v$RM_11863_out0 = v$S_9423_out0;
assign v$G1_7814_out0 = ((v$RD_5959_out0 && !v$RM_11399_out0) || (!v$RD_5959_out0) && v$RM_11399_out0);
assign v$G1_8278_out0 = ((v$RD_6423_out0 && !v$RM_11863_out0) || (!v$RD_6423_out0) && v$RM_11863_out0);
assign v$G2_12350_out0 = v$RD_5959_out0 && v$RM_11399_out0;
assign v$G2_12814_out0 = v$RD_6423_out0 && v$RM_11863_out0;
assign v$CARRY_4959_out0 = v$G2_12350_out0;
assign v$CARRY_5423_out0 = v$G2_12814_out0;
assign v$S_8960_out0 = v$G1_7814_out0;
assign v$S_9424_out0 = v$G1_8278_out0;
assign v$S_1265_out0 = v$S_8960_out0;
assign v$S_1489_out0 = v$S_9424_out0;
assign v$G1_4041_out0 = v$CARRY_4959_out0 || v$CARRY_4958_out0;
assign v$G1_4265_out0 = v$CARRY_5423_out0 || v$CARRY_5422_out0;
assign v$COUT_733_out0 = v$G1_4041_out0;
assign v$COUT_957_out0 = v$G1_4265_out0;
assign v$_10654_out0 = { v$_4552_out0,v$S_1265_out0 };
assign v$_10669_out0 = { v$_4567_out0,v$S_1489_out0 };
assign v$_10949_out0 = { v$_10654_out0,v$COUT_733_out0 };
assign v$_10964_out0 = { v$_10669_out0,v$COUT_957_out0 };
assign v$COUT_10919_out0 = v$_10949_out0;
assign v$COUT_10934_out0 = v$_10964_out0;
assign v$CIN_2363_out0 = v$COUT_10919_out0;
assign v$CIN_2378_out0 = v$COUT_10934_out0;
assign v$_476_out0 = v$CIN_2363_out0[8:8];
assign v$_491_out0 = v$CIN_2378_out0[8:8];
assign v$_1781_out0 = v$CIN_2363_out0[6:6];
assign v$_1796_out0 = v$CIN_2378_out0[6:6];
assign v$_2163_out0 = v$CIN_2363_out0[3:3];
assign v$_2178_out0 = v$CIN_2378_out0[3:3];
assign v$_2202_out0 = v$CIN_2363_out0[15:15];
assign v$_2216_out0 = v$CIN_2378_out0[15:15];
assign v$_2510_out0 = v$CIN_2363_out0[0:0];
assign v$_2525_out0 = v$CIN_2378_out0[0:0];
assign v$_3059_out0 = v$CIN_2363_out0[9:9];
assign v$_3074_out0 = v$CIN_2378_out0[9:9];
assign v$_3093_out0 = v$CIN_2363_out0[2:2];
assign v$_3108_out0 = v$CIN_2378_out0[2:2];
assign v$_3147_out0 = v$CIN_2363_out0[7:7];
assign v$_3162_out0 = v$CIN_2378_out0[7:7];
assign v$_3831_out0 = v$CIN_2363_out0[1:1];
assign v$_3846_out0 = v$CIN_2378_out0[1:1];
assign v$_3869_out0 = v$CIN_2363_out0[10:10];
assign v$_3884_out0 = v$CIN_2378_out0[10:10];
assign v$_6808_out0 = v$CIN_2363_out0[11:11];
assign v$_6823_out0 = v$CIN_2378_out0[11:11];
assign v$_7652_out0 = v$CIN_2363_out0[12:12];
assign v$_7667_out0 = v$CIN_2378_out0[12:12];
assign v$_8707_out0 = v$CIN_2363_out0[13:13];
assign v$_8722_out0 = v$CIN_2378_out0[13:13];
assign v$_8777_out0 = v$CIN_2363_out0[14:14];
assign v$_8792_out0 = v$CIN_2378_out0[14:14];
assign v$_10727_out0 = v$CIN_2363_out0[5:5];
assign v$_10742_out0 = v$CIN_2378_out0[5:5];
assign v$_13456_out0 = v$CIN_2363_out0[4:4];
assign v$_13471_out0 = v$CIN_2378_out0[4:4];
assign v$RM_3474_out0 = v$_7652_out0;
assign v$RM_3475_out0 = v$_8777_out0;
assign v$RM_3477_out0 = v$_10727_out0;
assign v$RM_3478_out0 = v$_13456_out0;
assign v$RM_3479_out0 = v$_8707_out0;
assign v$RM_3480_out0 = v$_3059_out0;
assign v$RM_3481_out0 = v$_3869_out0;
assign v$RM_3482_out0 = v$_3831_out0;
assign v$RM_3483_out0 = v$_2163_out0;
assign v$RM_3484_out0 = v$_1781_out0;
assign v$RM_3485_out0 = v$_3147_out0;
assign v$RM_3486_out0 = v$_6808_out0;
assign v$RM_3487_out0 = v$_476_out0;
assign v$RM_3488_out0 = v$_3093_out0;
assign v$RM_3698_out0 = v$_7667_out0;
assign v$RM_3699_out0 = v$_8792_out0;
assign v$RM_3701_out0 = v$_10742_out0;
assign v$RM_3702_out0 = v$_13471_out0;
assign v$RM_3703_out0 = v$_8722_out0;
assign v$RM_3704_out0 = v$_3074_out0;
assign v$RM_3705_out0 = v$_3884_out0;
assign v$RM_3706_out0 = v$_3846_out0;
assign v$RM_3707_out0 = v$_2178_out0;
assign v$RM_3708_out0 = v$_1796_out0;
assign v$RM_3709_out0 = v$_3162_out0;
assign v$RM_3710_out0 = v$_6823_out0;
assign v$RM_3711_out0 = v$_491_out0;
assign v$RM_3712_out0 = v$_3108_out0;
assign v$CIN_9929_out0 = v$_2202_out0;
assign v$CIN_10153_out0 = v$_2216_out0;
assign v$RM_11561_out0 = v$_2510_out0;
assign v$RM_12025_out0 = v$_2525_out0;
assign v$RD_6114_out0 = v$CIN_9929_out0;
assign v$RD_6578_out0 = v$CIN_10153_out0;
assign v$G1_7976_out0 = ((v$RD_6121_out0 && !v$RM_11561_out0) || (!v$RD_6121_out0) && v$RM_11561_out0);
assign v$G1_8440_out0 = ((v$RD_6585_out0 && !v$RM_12025_out0) || (!v$RD_6585_out0) && v$RM_12025_out0);
assign v$RM_11549_out0 = v$RM_3474_out0;
assign v$RM_11551_out0 = v$RM_3475_out0;
assign v$RM_11555_out0 = v$RM_3477_out0;
assign v$RM_11557_out0 = v$RM_3478_out0;
assign v$RM_11559_out0 = v$RM_3479_out0;
assign v$RM_11562_out0 = v$RM_3480_out0;
assign v$RM_11564_out0 = v$RM_3481_out0;
assign v$RM_11566_out0 = v$RM_3482_out0;
assign v$RM_11568_out0 = v$RM_3483_out0;
assign v$RM_11570_out0 = v$RM_3484_out0;
assign v$RM_11572_out0 = v$RM_3485_out0;
assign v$RM_11574_out0 = v$RM_3486_out0;
assign v$RM_11576_out0 = v$RM_3487_out0;
assign v$RM_11578_out0 = v$RM_3488_out0;
assign v$RM_12013_out0 = v$RM_3698_out0;
assign v$RM_12015_out0 = v$RM_3699_out0;
assign v$RM_12019_out0 = v$RM_3701_out0;
assign v$RM_12021_out0 = v$RM_3702_out0;
assign v$RM_12023_out0 = v$RM_3703_out0;
assign v$RM_12026_out0 = v$RM_3704_out0;
assign v$RM_12028_out0 = v$RM_3705_out0;
assign v$RM_12030_out0 = v$RM_3706_out0;
assign v$RM_12032_out0 = v$RM_3707_out0;
assign v$RM_12034_out0 = v$RM_3708_out0;
assign v$RM_12036_out0 = v$RM_3709_out0;
assign v$RM_12038_out0 = v$RM_3710_out0;
assign v$RM_12040_out0 = v$RM_3711_out0;
assign v$RM_12042_out0 = v$RM_3712_out0;
assign v$G2_12512_out0 = v$RD_6121_out0 && v$RM_11561_out0;
assign v$G2_12976_out0 = v$RD_6585_out0 && v$RM_12025_out0;
assign v$CARRY_5121_out0 = v$G2_12512_out0;
assign v$CARRY_5585_out0 = v$G2_12976_out0;
assign v$G1_7964_out0 = ((v$RD_6109_out0 && !v$RM_11549_out0) || (!v$RD_6109_out0) && v$RM_11549_out0);
assign v$G1_7966_out0 = ((v$RD_6111_out0 && !v$RM_11551_out0) || (!v$RD_6111_out0) && v$RM_11551_out0);
assign v$G1_7970_out0 = ((v$RD_6115_out0 && !v$RM_11555_out0) || (!v$RD_6115_out0) && v$RM_11555_out0);
assign v$G1_7972_out0 = ((v$RD_6117_out0 && !v$RM_11557_out0) || (!v$RD_6117_out0) && v$RM_11557_out0);
assign v$G1_7974_out0 = ((v$RD_6119_out0 && !v$RM_11559_out0) || (!v$RD_6119_out0) && v$RM_11559_out0);
assign v$G1_7977_out0 = ((v$RD_6122_out0 && !v$RM_11562_out0) || (!v$RD_6122_out0) && v$RM_11562_out0);
assign v$G1_7979_out0 = ((v$RD_6124_out0 && !v$RM_11564_out0) || (!v$RD_6124_out0) && v$RM_11564_out0);
assign v$G1_7981_out0 = ((v$RD_6126_out0 && !v$RM_11566_out0) || (!v$RD_6126_out0) && v$RM_11566_out0);
assign v$G1_7983_out0 = ((v$RD_6128_out0 && !v$RM_11568_out0) || (!v$RD_6128_out0) && v$RM_11568_out0);
assign v$G1_7985_out0 = ((v$RD_6130_out0 && !v$RM_11570_out0) || (!v$RD_6130_out0) && v$RM_11570_out0);
assign v$G1_7987_out0 = ((v$RD_6132_out0 && !v$RM_11572_out0) || (!v$RD_6132_out0) && v$RM_11572_out0);
assign v$G1_7989_out0 = ((v$RD_6134_out0 && !v$RM_11574_out0) || (!v$RD_6134_out0) && v$RM_11574_out0);
assign v$G1_7991_out0 = ((v$RD_6136_out0 && !v$RM_11576_out0) || (!v$RD_6136_out0) && v$RM_11576_out0);
assign v$G1_7993_out0 = ((v$RD_6138_out0 && !v$RM_11578_out0) || (!v$RD_6138_out0) && v$RM_11578_out0);
assign v$G1_8428_out0 = ((v$RD_6573_out0 && !v$RM_12013_out0) || (!v$RD_6573_out0) && v$RM_12013_out0);
assign v$G1_8430_out0 = ((v$RD_6575_out0 && !v$RM_12015_out0) || (!v$RD_6575_out0) && v$RM_12015_out0);
assign v$G1_8434_out0 = ((v$RD_6579_out0 && !v$RM_12019_out0) || (!v$RD_6579_out0) && v$RM_12019_out0);
assign v$G1_8436_out0 = ((v$RD_6581_out0 && !v$RM_12021_out0) || (!v$RD_6581_out0) && v$RM_12021_out0);
assign v$G1_8438_out0 = ((v$RD_6583_out0 && !v$RM_12023_out0) || (!v$RD_6583_out0) && v$RM_12023_out0);
assign v$G1_8441_out0 = ((v$RD_6586_out0 && !v$RM_12026_out0) || (!v$RD_6586_out0) && v$RM_12026_out0);
assign v$G1_8443_out0 = ((v$RD_6588_out0 && !v$RM_12028_out0) || (!v$RD_6588_out0) && v$RM_12028_out0);
assign v$G1_8445_out0 = ((v$RD_6590_out0 && !v$RM_12030_out0) || (!v$RD_6590_out0) && v$RM_12030_out0);
assign v$G1_8447_out0 = ((v$RD_6592_out0 && !v$RM_12032_out0) || (!v$RD_6592_out0) && v$RM_12032_out0);
assign v$G1_8449_out0 = ((v$RD_6594_out0 && !v$RM_12034_out0) || (!v$RD_6594_out0) && v$RM_12034_out0);
assign v$G1_8451_out0 = ((v$RD_6596_out0 && !v$RM_12036_out0) || (!v$RD_6596_out0) && v$RM_12036_out0);
assign v$G1_8453_out0 = ((v$RD_6598_out0 && !v$RM_12038_out0) || (!v$RD_6598_out0) && v$RM_12038_out0);
assign v$G1_8455_out0 = ((v$RD_6600_out0 && !v$RM_12040_out0) || (!v$RD_6600_out0) && v$RM_12040_out0);
assign v$G1_8457_out0 = ((v$RD_6602_out0 && !v$RM_12042_out0) || (!v$RD_6602_out0) && v$RM_12042_out0);
assign v$S_9122_out0 = v$G1_7976_out0;
assign v$S_9586_out0 = v$G1_8440_out0;
assign v$G2_12500_out0 = v$RD_6109_out0 && v$RM_11549_out0;
assign v$G2_12502_out0 = v$RD_6111_out0 && v$RM_11551_out0;
assign v$G2_12506_out0 = v$RD_6115_out0 && v$RM_11555_out0;
assign v$G2_12508_out0 = v$RD_6117_out0 && v$RM_11557_out0;
assign v$G2_12510_out0 = v$RD_6119_out0 && v$RM_11559_out0;
assign v$G2_12513_out0 = v$RD_6122_out0 && v$RM_11562_out0;
assign v$G2_12515_out0 = v$RD_6124_out0 && v$RM_11564_out0;
assign v$G2_12517_out0 = v$RD_6126_out0 && v$RM_11566_out0;
assign v$G2_12519_out0 = v$RD_6128_out0 && v$RM_11568_out0;
assign v$G2_12521_out0 = v$RD_6130_out0 && v$RM_11570_out0;
assign v$G2_12523_out0 = v$RD_6132_out0 && v$RM_11572_out0;
assign v$G2_12525_out0 = v$RD_6134_out0 && v$RM_11574_out0;
assign v$G2_12527_out0 = v$RD_6136_out0 && v$RM_11576_out0;
assign v$G2_12529_out0 = v$RD_6138_out0 && v$RM_11578_out0;
assign v$G2_12964_out0 = v$RD_6573_out0 && v$RM_12013_out0;
assign v$G2_12966_out0 = v$RD_6575_out0 && v$RM_12015_out0;
assign v$G2_12970_out0 = v$RD_6579_out0 && v$RM_12019_out0;
assign v$G2_12972_out0 = v$RD_6581_out0 && v$RM_12021_out0;
assign v$G2_12974_out0 = v$RD_6583_out0 && v$RM_12023_out0;
assign v$G2_12977_out0 = v$RD_6586_out0 && v$RM_12026_out0;
assign v$G2_12979_out0 = v$RD_6588_out0 && v$RM_12028_out0;
assign v$G2_12981_out0 = v$RD_6590_out0 && v$RM_12030_out0;
assign v$G2_12983_out0 = v$RD_6592_out0 && v$RM_12032_out0;
assign v$G2_12985_out0 = v$RD_6594_out0 && v$RM_12034_out0;
assign v$G2_12987_out0 = v$RD_6596_out0 && v$RM_12036_out0;
assign v$G2_12989_out0 = v$RD_6598_out0 && v$RM_12038_out0;
assign v$G2_12991_out0 = v$RD_6600_out0 && v$RM_12040_out0;
assign v$G2_12993_out0 = v$RD_6602_out0 && v$RM_12042_out0;
assign v$S_4673_out0 = v$S_9122_out0;
assign v$S_4688_out0 = v$S_9586_out0;
assign v$CARRY_5109_out0 = v$G2_12500_out0;
assign v$CARRY_5111_out0 = v$G2_12502_out0;
assign v$CARRY_5115_out0 = v$G2_12506_out0;
assign v$CARRY_5117_out0 = v$G2_12508_out0;
assign v$CARRY_5119_out0 = v$G2_12510_out0;
assign v$CARRY_5122_out0 = v$G2_12513_out0;
assign v$CARRY_5124_out0 = v$G2_12515_out0;
assign v$CARRY_5126_out0 = v$G2_12517_out0;
assign v$CARRY_5128_out0 = v$G2_12519_out0;
assign v$CARRY_5130_out0 = v$G2_12521_out0;
assign v$CARRY_5132_out0 = v$G2_12523_out0;
assign v$CARRY_5134_out0 = v$G2_12525_out0;
assign v$CARRY_5136_out0 = v$G2_12527_out0;
assign v$CARRY_5138_out0 = v$G2_12529_out0;
assign v$CARRY_5573_out0 = v$G2_12964_out0;
assign v$CARRY_5575_out0 = v$G2_12966_out0;
assign v$CARRY_5579_out0 = v$G2_12970_out0;
assign v$CARRY_5581_out0 = v$G2_12972_out0;
assign v$CARRY_5583_out0 = v$G2_12974_out0;
assign v$CARRY_5586_out0 = v$G2_12977_out0;
assign v$CARRY_5588_out0 = v$G2_12979_out0;
assign v$CARRY_5590_out0 = v$G2_12981_out0;
assign v$CARRY_5592_out0 = v$G2_12983_out0;
assign v$CARRY_5594_out0 = v$G2_12985_out0;
assign v$CARRY_5596_out0 = v$G2_12987_out0;
assign v$CARRY_5598_out0 = v$G2_12989_out0;
assign v$CARRY_5600_out0 = v$G2_12991_out0;
assign v$CARRY_5602_out0 = v$G2_12993_out0;
assign v$S_9110_out0 = v$G1_7964_out0;
assign v$S_9112_out0 = v$G1_7966_out0;
assign v$S_9116_out0 = v$G1_7970_out0;
assign v$S_9118_out0 = v$G1_7972_out0;
assign v$S_9120_out0 = v$G1_7974_out0;
assign v$S_9123_out0 = v$G1_7977_out0;
assign v$S_9125_out0 = v$G1_7979_out0;
assign v$S_9127_out0 = v$G1_7981_out0;
assign v$S_9129_out0 = v$G1_7983_out0;
assign v$S_9131_out0 = v$G1_7985_out0;
assign v$S_9133_out0 = v$G1_7987_out0;
assign v$S_9135_out0 = v$G1_7989_out0;
assign v$S_9137_out0 = v$G1_7991_out0;
assign v$S_9139_out0 = v$G1_7993_out0;
assign v$S_9574_out0 = v$G1_8428_out0;
assign v$S_9576_out0 = v$G1_8430_out0;
assign v$S_9580_out0 = v$G1_8434_out0;
assign v$S_9582_out0 = v$G1_8436_out0;
assign v$S_9584_out0 = v$G1_8438_out0;
assign v$S_9587_out0 = v$G1_8441_out0;
assign v$S_9589_out0 = v$G1_8443_out0;
assign v$S_9591_out0 = v$G1_8445_out0;
assign v$S_9593_out0 = v$G1_8447_out0;
assign v$S_9595_out0 = v$G1_8449_out0;
assign v$S_9597_out0 = v$G1_8451_out0;
assign v$S_9599_out0 = v$G1_8453_out0;
assign v$S_9601_out0 = v$G1_8455_out0;
assign v$S_9603_out0 = v$G1_8457_out0;
assign v$CIN_9935_out0 = v$CARRY_5121_out0;
assign v$CIN_10159_out0 = v$CARRY_5585_out0;
assign v$RD_6127_out0 = v$CIN_9935_out0;
assign v$RD_6591_out0 = v$CIN_10159_out0;
assign v$_9802_out0 = { v$_2439_out0,v$S_4673_out0 };
assign v$_9803_out0 = { v$_2440_out0,v$S_4688_out0 };
assign v$RM_11550_out0 = v$S_9110_out0;
assign v$RM_11552_out0 = v$S_9112_out0;
assign v$RM_11556_out0 = v$S_9116_out0;
assign v$RM_11558_out0 = v$S_9118_out0;
assign v$RM_11560_out0 = v$S_9120_out0;
assign v$RM_11563_out0 = v$S_9123_out0;
assign v$RM_11565_out0 = v$S_9125_out0;
assign v$RM_11567_out0 = v$S_9127_out0;
assign v$RM_11569_out0 = v$S_9129_out0;
assign v$RM_11571_out0 = v$S_9131_out0;
assign v$RM_11573_out0 = v$S_9133_out0;
assign v$RM_11575_out0 = v$S_9135_out0;
assign v$RM_11577_out0 = v$S_9137_out0;
assign v$RM_11579_out0 = v$S_9139_out0;
assign v$RM_12014_out0 = v$S_9574_out0;
assign v$RM_12016_out0 = v$S_9576_out0;
assign v$RM_12020_out0 = v$S_9580_out0;
assign v$RM_12022_out0 = v$S_9582_out0;
assign v$RM_12024_out0 = v$S_9584_out0;
assign v$RM_12027_out0 = v$S_9587_out0;
assign v$RM_12029_out0 = v$S_9589_out0;
assign v$RM_12031_out0 = v$S_9591_out0;
assign v$RM_12033_out0 = v$S_9593_out0;
assign v$RM_12035_out0 = v$S_9595_out0;
assign v$RM_12037_out0 = v$S_9597_out0;
assign v$RM_12039_out0 = v$S_9599_out0;
assign v$RM_12041_out0 = v$S_9601_out0;
assign v$RM_12043_out0 = v$S_9603_out0;
assign v$G1_7982_out0 = ((v$RD_6127_out0 && !v$RM_11567_out0) || (!v$RD_6127_out0) && v$RM_11567_out0);
assign v$G1_8446_out0 = ((v$RD_6591_out0 && !v$RM_12031_out0) || (!v$RD_6591_out0) && v$RM_12031_out0);
assign v$G2_12518_out0 = v$RD_6127_out0 && v$RM_11567_out0;
assign v$G2_12982_out0 = v$RD_6591_out0 && v$RM_12031_out0;
assign v$CARRY_5127_out0 = v$G2_12518_out0;
assign v$CARRY_5591_out0 = v$G2_12982_out0;
assign v$S_9128_out0 = v$G1_7982_out0;
assign v$S_9592_out0 = v$G1_8446_out0;
assign v$S_1346_out0 = v$S_9128_out0;
assign v$S_1570_out0 = v$S_9592_out0;
assign v$G1_4122_out0 = v$CARRY_5127_out0 || v$CARRY_5126_out0;
assign v$G1_4346_out0 = v$CARRY_5591_out0 || v$CARRY_5590_out0;
assign v$COUT_814_out0 = v$G1_4122_out0;
assign v$COUT_1038_out0 = v$G1_4346_out0;
assign v$CIN_9941_out0 = v$COUT_814_out0;
assign v$CIN_10165_out0 = v$COUT_1038_out0;
assign v$RD_6139_out0 = v$CIN_9941_out0;
assign v$RD_6603_out0 = v$CIN_10165_out0;
assign v$G1_7994_out0 = ((v$RD_6139_out0 && !v$RM_11579_out0) || (!v$RD_6139_out0) && v$RM_11579_out0);
assign v$G1_8458_out0 = ((v$RD_6603_out0 && !v$RM_12043_out0) || (!v$RD_6603_out0) && v$RM_12043_out0);
assign v$G2_12530_out0 = v$RD_6139_out0 && v$RM_11579_out0;
assign v$G2_12994_out0 = v$RD_6603_out0 && v$RM_12043_out0;
assign v$CARRY_5139_out0 = v$G2_12530_out0;
assign v$CARRY_5603_out0 = v$G2_12994_out0;
assign v$S_9140_out0 = v$G1_7994_out0;
assign v$S_9604_out0 = v$G1_8458_out0;
assign v$S_1352_out0 = v$S_9140_out0;
assign v$S_1576_out0 = v$S_9604_out0;
assign v$G1_4128_out0 = v$CARRY_5139_out0 || v$CARRY_5138_out0;
assign v$G1_4352_out0 = v$CARRY_5603_out0 || v$CARRY_5602_out0;
assign v$COUT_820_out0 = v$G1_4128_out0;
assign v$COUT_1044_out0 = v$G1_4352_out0;
assign v$_4790_out0 = { v$S_1346_out0,v$S_1352_out0 };
assign v$_4805_out0 = { v$S_1570_out0,v$S_1576_out0 };
assign v$CIN_9936_out0 = v$COUT_820_out0;
assign v$CIN_10160_out0 = v$COUT_1044_out0;
assign v$RD_6129_out0 = v$CIN_9936_out0;
assign v$RD_6593_out0 = v$CIN_10160_out0;
assign v$G1_7984_out0 = ((v$RD_6129_out0 && !v$RM_11569_out0) || (!v$RD_6129_out0) && v$RM_11569_out0);
assign v$G1_8448_out0 = ((v$RD_6593_out0 && !v$RM_12033_out0) || (!v$RD_6593_out0) && v$RM_12033_out0);
assign v$G2_12520_out0 = v$RD_6129_out0 && v$RM_11569_out0;
assign v$G2_12984_out0 = v$RD_6593_out0 && v$RM_12033_out0;
assign v$CARRY_5129_out0 = v$G2_12520_out0;
assign v$CARRY_5593_out0 = v$G2_12984_out0;
assign v$S_9130_out0 = v$G1_7984_out0;
assign v$S_9594_out0 = v$G1_8448_out0;
assign v$S_1347_out0 = v$S_9130_out0;
assign v$S_1571_out0 = v$S_9594_out0;
assign v$G1_4123_out0 = v$CARRY_5129_out0 || v$CARRY_5128_out0;
assign v$G1_4347_out0 = v$CARRY_5593_out0 || v$CARRY_5592_out0;
assign v$COUT_815_out0 = v$G1_4123_out0;
assign v$COUT_1039_out0 = v$G1_4347_out0;
assign v$_2560_out0 = { v$_4790_out0,v$S_1347_out0 };
assign v$_2575_out0 = { v$_4805_out0,v$S_1571_out0 };
assign v$CIN_9931_out0 = v$COUT_815_out0;
assign v$CIN_10155_out0 = v$COUT_1039_out0;
assign v$RD_6118_out0 = v$CIN_9931_out0;
assign v$RD_6582_out0 = v$CIN_10155_out0;
assign v$G1_7973_out0 = ((v$RD_6118_out0 && !v$RM_11558_out0) || (!v$RD_6118_out0) && v$RM_11558_out0);
assign v$G1_8437_out0 = ((v$RD_6582_out0 && !v$RM_12022_out0) || (!v$RD_6582_out0) && v$RM_12022_out0);
assign v$G2_12509_out0 = v$RD_6118_out0 && v$RM_11558_out0;
assign v$G2_12973_out0 = v$RD_6582_out0 && v$RM_12022_out0;
assign v$CARRY_5118_out0 = v$G2_12509_out0;
assign v$CARRY_5582_out0 = v$G2_12973_out0;
assign v$S_9119_out0 = v$G1_7973_out0;
assign v$S_9583_out0 = v$G1_8437_out0;
assign v$S_1342_out0 = v$S_9119_out0;
assign v$S_1566_out0 = v$S_9583_out0;
assign v$G1_4118_out0 = v$CARRY_5118_out0 || v$CARRY_5117_out0;
assign v$G1_4342_out0 = v$CARRY_5582_out0 || v$CARRY_5581_out0;
assign v$COUT_810_out0 = v$G1_4118_out0;
assign v$COUT_1034_out0 = v$G1_4342_out0;
assign v$_7040_out0 = { v$_2560_out0,v$S_1342_out0 };
assign v$_7055_out0 = { v$_2575_out0,v$S_1566_out0 };
assign v$CIN_9930_out0 = v$COUT_810_out0;
assign v$CIN_10154_out0 = v$COUT_1034_out0;
assign v$RD_6116_out0 = v$CIN_9930_out0;
assign v$RD_6580_out0 = v$CIN_10154_out0;
assign v$G1_7971_out0 = ((v$RD_6116_out0 && !v$RM_11556_out0) || (!v$RD_6116_out0) && v$RM_11556_out0);
assign v$G1_8435_out0 = ((v$RD_6580_out0 && !v$RM_12020_out0) || (!v$RD_6580_out0) && v$RM_12020_out0);
assign v$G2_12507_out0 = v$RD_6116_out0 && v$RM_11556_out0;
assign v$G2_12971_out0 = v$RD_6580_out0 && v$RM_12020_out0;
assign v$CARRY_5116_out0 = v$G2_12507_out0;
assign v$CARRY_5580_out0 = v$G2_12971_out0;
assign v$S_9117_out0 = v$G1_7971_out0;
assign v$S_9581_out0 = v$G1_8435_out0;
assign v$S_1341_out0 = v$S_9117_out0;
assign v$S_1565_out0 = v$S_9581_out0;
assign v$G1_4117_out0 = v$CARRY_5116_out0 || v$CARRY_5115_out0;
assign v$G1_4341_out0 = v$CARRY_5580_out0 || v$CARRY_5579_out0;
assign v$COUT_809_out0 = v$G1_4117_out0;
assign v$COUT_1033_out0 = v$G1_4341_out0;
assign v$_13526_out0 = { v$_7040_out0,v$S_1341_out0 };
assign v$_13541_out0 = { v$_7055_out0,v$S_1565_out0 };
assign v$CIN_9937_out0 = v$COUT_809_out0;
assign v$CIN_10161_out0 = v$COUT_1033_out0;
assign v$RD_6131_out0 = v$CIN_9937_out0;
assign v$RD_6595_out0 = v$CIN_10161_out0;
assign v$G1_7986_out0 = ((v$RD_6131_out0 && !v$RM_11571_out0) || (!v$RD_6131_out0) && v$RM_11571_out0);
assign v$G1_8450_out0 = ((v$RD_6595_out0 && !v$RM_12035_out0) || (!v$RD_6595_out0) && v$RM_12035_out0);
assign v$G2_12522_out0 = v$RD_6131_out0 && v$RM_11571_out0;
assign v$G2_12986_out0 = v$RD_6595_out0 && v$RM_12035_out0;
assign v$CARRY_5131_out0 = v$G2_12522_out0;
assign v$CARRY_5595_out0 = v$G2_12986_out0;
assign v$S_9132_out0 = v$G1_7986_out0;
assign v$S_9596_out0 = v$G1_8450_out0;
assign v$S_1348_out0 = v$S_9132_out0;
assign v$S_1572_out0 = v$S_9596_out0;
assign v$G1_4124_out0 = v$CARRY_5131_out0 || v$CARRY_5130_out0;
assign v$G1_4348_out0 = v$CARRY_5595_out0 || v$CARRY_5594_out0;
assign v$COUT_816_out0 = v$G1_4124_out0;
assign v$COUT_1040_out0 = v$G1_4348_out0;
assign v$_3319_out0 = { v$_13526_out0,v$S_1348_out0 };
assign v$_3334_out0 = { v$_13541_out0,v$S_1572_out0 };
assign v$CIN_9938_out0 = v$COUT_816_out0;
assign v$CIN_10162_out0 = v$COUT_1040_out0;
assign v$RD_6133_out0 = v$CIN_9938_out0;
assign v$RD_6597_out0 = v$CIN_10162_out0;
assign v$G1_7988_out0 = ((v$RD_6133_out0 && !v$RM_11573_out0) || (!v$RD_6133_out0) && v$RM_11573_out0);
assign v$G1_8452_out0 = ((v$RD_6597_out0 && !v$RM_12037_out0) || (!v$RD_6597_out0) && v$RM_12037_out0);
assign v$G2_12524_out0 = v$RD_6133_out0 && v$RM_11573_out0;
assign v$G2_12988_out0 = v$RD_6597_out0 && v$RM_12037_out0;
assign v$CARRY_5133_out0 = v$G2_12524_out0;
assign v$CARRY_5597_out0 = v$G2_12988_out0;
assign v$S_9134_out0 = v$G1_7988_out0;
assign v$S_9598_out0 = v$G1_8452_out0;
assign v$S_1349_out0 = v$S_9134_out0;
assign v$S_1573_out0 = v$S_9598_out0;
assign v$G1_4125_out0 = v$CARRY_5133_out0 || v$CARRY_5132_out0;
assign v$G1_4349_out0 = v$CARRY_5597_out0 || v$CARRY_5596_out0;
assign v$COUT_817_out0 = v$G1_4125_out0;
assign v$COUT_1041_out0 = v$G1_4349_out0;
assign v$_7155_out0 = { v$_3319_out0,v$S_1349_out0 };
assign v$_7170_out0 = { v$_3334_out0,v$S_1573_out0 };
assign v$CIN_9940_out0 = v$COUT_817_out0;
assign v$CIN_10164_out0 = v$COUT_1041_out0;
assign v$RD_6137_out0 = v$CIN_9940_out0;
assign v$RD_6601_out0 = v$CIN_10164_out0;
assign v$G1_7992_out0 = ((v$RD_6137_out0 && !v$RM_11577_out0) || (!v$RD_6137_out0) && v$RM_11577_out0);
assign v$G1_8456_out0 = ((v$RD_6601_out0 && !v$RM_12041_out0) || (!v$RD_6601_out0) && v$RM_12041_out0);
assign v$G2_12528_out0 = v$RD_6137_out0 && v$RM_11577_out0;
assign v$G2_12992_out0 = v$RD_6601_out0 && v$RM_12041_out0;
assign v$CARRY_5137_out0 = v$G2_12528_out0;
assign v$CARRY_5601_out0 = v$G2_12992_out0;
assign v$S_9138_out0 = v$G1_7992_out0;
assign v$S_9602_out0 = v$G1_8456_out0;
assign v$S_1351_out0 = v$S_9138_out0;
assign v$S_1575_out0 = v$S_9602_out0;
assign v$G1_4127_out0 = v$CARRY_5137_out0 || v$CARRY_5136_out0;
assign v$G1_4351_out0 = v$CARRY_5601_out0 || v$CARRY_5600_out0;
assign v$COUT_819_out0 = v$G1_4127_out0;
assign v$COUT_1043_out0 = v$G1_4351_out0;
assign v$_4757_out0 = { v$_7155_out0,v$S_1351_out0 };
assign v$_4772_out0 = { v$_7170_out0,v$S_1575_out0 };
assign v$CIN_9933_out0 = v$COUT_819_out0;
assign v$CIN_10157_out0 = v$COUT_1043_out0;
assign v$RD_6123_out0 = v$CIN_9933_out0;
assign v$RD_6587_out0 = v$CIN_10157_out0;
assign v$G1_7978_out0 = ((v$RD_6123_out0 && !v$RM_11563_out0) || (!v$RD_6123_out0) && v$RM_11563_out0);
assign v$G1_8442_out0 = ((v$RD_6587_out0 && !v$RM_12027_out0) || (!v$RD_6587_out0) && v$RM_12027_out0);
assign v$G2_12514_out0 = v$RD_6123_out0 && v$RM_11563_out0;
assign v$G2_12978_out0 = v$RD_6587_out0 && v$RM_12027_out0;
assign v$CARRY_5123_out0 = v$G2_12514_out0;
assign v$CARRY_5587_out0 = v$G2_12978_out0;
assign v$S_9124_out0 = v$G1_7978_out0;
assign v$S_9588_out0 = v$G1_8442_out0;
assign v$S_1344_out0 = v$S_9124_out0;
assign v$S_1568_out0 = v$S_9588_out0;
assign v$G1_4120_out0 = v$CARRY_5123_out0 || v$CARRY_5122_out0;
assign v$G1_4344_out0 = v$CARRY_5587_out0 || v$CARRY_5586_out0;
assign v$COUT_812_out0 = v$G1_4120_out0;
assign v$COUT_1036_out0 = v$G1_4344_out0;
assign v$_6934_out0 = { v$_4757_out0,v$S_1344_out0 };
assign v$_6949_out0 = { v$_4772_out0,v$S_1568_out0 };
assign v$CIN_9934_out0 = v$COUT_812_out0;
assign v$CIN_10158_out0 = v$COUT_1036_out0;
assign v$RD_6125_out0 = v$CIN_9934_out0;
assign v$RD_6589_out0 = v$CIN_10158_out0;
assign v$G1_7980_out0 = ((v$RD_6125_out0 && !v$RM_11565_out0) || (!v$RD_6125_out0) && v$RM_11565_out0);
assign v$G1_8444_out0 = ((v$RD_6589_out0 && !v$RM_12029_out0) || (!v$RD_6589_out0) && v$RM_12029_out0);
assign v$G2_12516_out0 = v$RD_6125_out0 && v$RM_11565_out0;
assign v$G2_12980_out0 = v$RD_6589_out0 && v$RM_12029_out0;
assign v$CARRY_5125_out0 = v$G2_12516_out0;
assign v$CARRY_5589_out0 = v$G2_12980_out0;
assign v$S_9126_out0 = v$G1_7980_out0;
assign v$S_9590_out0 = v$G1_8444_out0;
assign v$S_1345_out0 = v$S_9126_out0;
assign v$S_1569_out0 = v$S_9590_out0;
assign v$G1_4121_out0 = v$CARRY_5125_out0 || v$CARRY_5124_out0;
assign v$G1_4345_out0 = v$CARRY_5589_out0 || v$CARRY_5588_out0;
assign v$COUT_813_out0 = v$G1_4121_out0;
assign v$COUT_1037_out0 = v$G1_4345_out0;
assign v$_5810_out0 = { v$_6934_out0,v$S_1345_out0 };
assign v$_5825_out0 = { v$_6949_out0,v$S_1569_out0 };
assign v$CIN_9939_out0 = v$COUT_813_out0;
assign v$CIN_10163_out0 = v$COUT_1037_out0;
assign v$RD_6135_out0 = v$CIN_9939_out0;
assign v$RD_6599_out0 = v$CIN_10163_out0;
assign v$G1_7990_out0 = ((v$RD_6135_out0 && !v$RM_11575_out0) || (!v$RD_6135_out0) && v$RM_11575_out0);
assign v$G1_8454_out0 = ((v$RD_6599_out0 && !v$RM_12039_out0) || (!v$RD_6599_out0) && v$RM_12039_out0);
assign v$G2_12526_out0 = v$RD_6135_out0 && v$RM_11575_out0;
assign v$G2_12990_out0 = v$RD_6599_out0 && v$RM_12039_out0;
assign v$CARRY_5135_out0 = v$G2_12526_out0;
assign v$CARRY_5599_out0 = v$G2_12990_out0;
assign v$S_9136_out0 = v$G1_7990_out0;
assign v$S_9600_out0 = v$G1_8454_out0;
assign v$S_1350_out0 = v$S_9136_out0;
assign v$S_1574_out0 = v$S_9600_out0;
assign v$G1_4126_out0 = v$CARRY_5135_out0 || v$CARRY_5134_out0;
assign v$G1_4350_out0 = v$CARRY_5599_out0 || v$CARRY_5598_out0;
assign v$COUT_818_out0 = v$G1_4126_out0;
assign v$COUT_1042_out0 = v$G1_4350_out0;
assign v$_2034_out0 = { v$_5810_out0,v$S_1350_out0 };
assign v$_2049_out0 = { v$_5825_out0,v$S_1574_out0 };
assign v$CIN_9927_out0 = v$COUT_818_out0;
assign v$CIN_10151_out0 = v$COUT_1042_out0;
assign v$RD_6110_out0 = v$CIN_9927_out0;
assign v$RD_6574_out0 = v$CIN_10151_out0;
assign v$G1_7965_out0 = ((v$RD_6110_out0 && !v$RM_11550_out0) || (!v$RD_6110_out0) && v$RM_11550_out0);
assign v$G1_8429_out0 = ((v$RD_6574_out0 && !v$RM_12014_out0) || (!v$RD_6574_out0) && v$RM_12014_out0);
assign v$G2_12501_out0 = v$RD_6110_out0 && v$RM_11550_out0;
assign v$G2_12965_out0 = v$RD_6574_out0 && v$RM_12014_out0;
assign v$CARRY_5110_out0 = v$G2_12501_out0;
assign v$CARRY_5574_out0 = v$G2_12965_out0;
assign v$S_9111_out0 = v$G1_7965_out0;
assign v$S_9575_out0 = v$G1_8429_out0;
assign v$S_1338_out0 = v$S_9111_out0;
assign v$S_1562_out0 = v$S_9575_out0;
assign v$G1_4114_out0 = v$CARRY_5110_out0 || v$CARRY_5109_out0;
assign v$G1_4338_out0 = v$CARRY_5574_out0 || v$CARRY_5573_out0;
assign v$COUT_806_out0 = v$G1_4114_out0;
assign v$COUT_1030_out0 = v$G1_4338_out0;
assign v$_2801_out0 = { v$_2034_out0,v$S_1338_out0 };
assign v$_2816_out0 = { v$_2049_out0,v$S_1562_out0 };
assign v$CIN_9932_out0 = v$COUT_806_out0;
assign v$CIN_10156_out0 = v$COUT_1030_out0;
assign v$RD_6120_out0 = v$CIN_9932_out0;
assign v$RD_6584_out0 = v$CIN_10156_out0;
assign v$G1_7975_out0 = ((v$RD_6120_out0 && !v$RM_11560_out0) || (!v$RD_6120_out0) && v$RM_11560_out0);
assign v$G1_8439_out0 = ((v$RD_6584_out0 && !v$RM_12024_out0) || (!v$RD_6584_out0) && v$RM_12024_out0);
assign v$G2_12511_out0 = v$RD_6120_out0 && v$RM_11560_out0;
assign v$G2_12975_out0 = v$RD_6584_out0 && v$RM_12024_out0;
assign v$CARRY_5120_out0 = v$G2_12511_out0;
assign v$CARRY_5584_out0 = v$G2_12975_out0;
assign v$S_9121_out0 = v$G1_7975_out0;
assign v$S_9585_out0 = v$G1_8439_out0;
assign v$S_1343_out0 = v$S_9121_out0;
assign v$S_1567_out0 = v$S_9585_out0;
assign v$G1_4119_out0 = v$CARRY_5120_out0 || v$CARRY_5119_out0;
assign v$G1_4343_out0 = v$CARRY_5584_out0 || v$CARRY_5583_out0;
assign v$COUT_811_out0 = v$G1_4119_out0;
assign v$COUT_1035_out0 = v$G1_4343_out0;
assign v$_1833_out0 = { v$_2801_out0,v$S_1343_out0 };
assign v$_1848_out0 = { v$_2816_out0,v$S_1567_out0 };
assign v$CIN_9928_out0 = v$COUT_811_out0;
assign v$CIN_10152_out0 = v$COUT_1035_out0;
assign v$RD_6112_out0 = v$CIN_9928_out0;
assign v$RD_6576_out0 = v$CIN_10152_out0;
assign v$G1_7967_out0 = ((v$RD_6112_out0 && !v$RM_11552_out0) || (!v$RD_6112_out0) && v$RM_11552_out0);
assign v$G1_8431_out0 = ((v$RD_6576_out0 && !v$RM_12016_out0) || (!v$RD_6576_out0) && v$RM_12016_out0);
assign v$G2_12503_out0 = v$RD_6112_out0 && v$RM_11552_out0;
assign v$G2_12967_out0 = v$RD_6576_out0 && v$RM_12016_out0;
assign v$CARRY_5112_out0 = v$G2_12503_out0;
assign v$CARRY_5576_out0 = v$G2_12967_out0;
assign v$S_9113_out0 = v$G1_7967_out0;
assign v$S_9577_out0 = v$G1_8431_out0;
assign v$S_1339_out0 = v$S_9113_out0;
assign v$S_1563_out0 = v$S_9577_out0;
assign v$G1_4115_out0 = v$CARRY_5112_out0 || v$CARRY_5111_out0;
assign v$G1_4339_out0 = v$CARRY_5576_out0 || v$CARRY_5575_out0;
assign v$COUT_807_out0 = v$G1_4115_out0;
assign v$COUT_1031_out0 = v$G1_4339_out0;
assign v$_4557_out0 = { v$_1833_out0,v$S_1339_out0 };
assign v$_4572_out0 = { v$_1848_out0,v$S_1563_out0 };
assign v$RM_3476_out0 = v$COUT_807_out0;
assign v$RM_3700_out0 = v$COUT_1031_out0;
assign v$RM_11553_out0 = v$RM_3476_out0;
assign v$RM_12017_out0 = v$RM_3700_out0;
assign v$G1_7968_out0 = ((v$RD_6113_out0 && !v$RM_11553_out0) || (!v$RD_6113_out0) && v$RM_11553_out0);
assign v$G1_8432_out0 = ((v$RD_6577_out0 && !v$RM_12017_out0) || (!v$RD_6577_out0) && v$RM_12017_out0);
assign v$G2_12504_out0 = v$RD_6113_out0 && v$RM_11553_out0;
assign v$G2_12968_out0 = v$RD_6577_out0 && v$RM_12017_out0;
assign v$CARRY_5113_out0 = v$G2_12504_out0;
assign v$CARRY_5577_out0 = v$G2_12968_out0;
assign v$S_9114_out0 = v$G1_7968_out0;
assign v$S_9578_out0 = v$G1_8432_out0;
assign v$RM_11554_out0 = v$S_9114_out0;
assign v$RM_12018_out0 = v$S_9578_out0;
assign v$G1_7969_out0 = ((v$RD_6114_out0 && !v$RM_11554_out0) || (!v$RD_6114_out0) && v$RM_11554_out0);
assign v$G1_8433_out0 = ((v$RD_6578_out0 && !v$RM_12018_out0) || (!v$RD_6578_out0) && v$RM_12018_out0);
assign v$G2_12505_out0 = v$RD_6114_out0 && v$RM_11554_out0;
assign v$G2_12969_out0 = v$RD_6578_out0 && v$RM_12018_out0;
assign v$CARRY_5114_out0 = v$G2_12505_out0;
assign v$CARRY_5578_out0 = v$G2_12969_out0;
assign v$S_9115_out0 = v$G1_7969_out0;
assign v$S_9579_out0 = v$G1_8433_out0;
assign v$S_1340_out0 = v$S_9115_out0;
assign v$S_1564_out0 = v$S_9579_out0;
assign v$G1_4116_out0 = v$CARRY_5114_out0 || v$CARRY_5113_out0;
assign v$G1_4340_out0 = v$CARRY_5578_out0 || v$CARRY_5577_out0;
assign v$COUT_808_out0 = v$G1_4116_out0;
assign v$COUT_1032_out0 = v$G1_4340_out0;
assign v$_10659_out0 = { v$_4557_out0,v$S_1340_out0 };
assign v$_10674_out0 = { v$_4572_out0,v$S_1564_out0 };
assign v$_10954_out0 = { v$_10659_out0,v$COUT_808_out0 };
assign v$_10969_out0 = { v$_10674_out0,v$COUT_1032_out0 };
assign v$COUT_10924_out0 = v$_10954_out0;
assign v$COUT_10939_out0 = v$_10969_out0;
assign v$CIN_2367_out0 = v$COUT_10924_out0;
assign v$CIN_2382_out0 = v$COUT_10939_out0;
assign v$_480_out0 = v$CIN_2367_out0[8:8];
assign v$_495_out0 = v$CIN_2382_out0[8:8];
assign v$_1785_out0 = v$CIN_2367_out0[6:6];
assign v$_1800_out0 = v$CIN_2382_out0[6:6];
assign v$_2167_out0 = v$CIN_2367_out0[3:3];
assign v$_2182_out0 = v$CIN_2382_out0[3:3];
assign v$_2206_out0 = v$CIN_2367_out0[15:15];
assign v$_2220_out0 = v$CIN_2382_out0[15:15];
assign v$_2514_out0 = v$CIN_2367_out0[0:0];
assign v$_2529_out0 = v$CIN_2382_out0[0:0];
assign v$_3063_out0 = v$CIN_2367_out0[9:9];
assign v$_3078_out0 = v$CIN_2382_out0[9:9];
assign v$_3097_out0 = v$CIN_2367_out0[2:2];
assign v$_3112_out0 = v$CIN_2382_out0[2:2];
assign v$_3151_out0 = v$CIN_2367_out0[7:7];
assign v$_3166_out0 = v$CIN_2382_out0[7:7];
assign v$_3835_out0 = v$CIN_2367_out0[1:1];
assign v$_3850_out0 = v$CIN_2382_out0[1:1];
assign v$_3873_out0 = v$CIN_2367_out0[10:10];
assign v$_3888_out0 = v$CIN_2382_out0[10:10];
assign v$_6812_out0 = v$CIN_2367_out0[11:11];
assign v$_6827_out0 = v$CIN_2382_out0[11:11];
assign v$_7656_out0 = v$CIN_2367_out0[12:12];
assign v$_7671_out0 = v$CIN_2382_out0[12:12];
assign v$_8711_out0 = v$CIN_2367_out0[13:13];
assign v$_8726_out0 = v$CIN_2382_out0[13:13];
assign v$_8781_out0 = v$CIN_2367_out0[14:14];
assign v$_8796_out0 = v$CIN_2382_out0[14:14];
assign v$_10731_out0 = v$CIN_2367_out0[5:5];
assign v$_10746_out0 = v$CIN_2382_out0[5:5];
assign v$_13460_out0 = v$CIN_2367_out0[4:4];
assign v$_13475_out0 = v$CIN_2382_out0[4:4];
assign v$RM_3534_out0 = v$_7656_out0;
assign v$RM_3535_out0 = v$_8781_out0;
assign v$RM_3537_out0 = v$_10731_out0;
assign v$RM_3538_out0 = v$_13460_out0;
assign v$RM_3539_out0 = v$_8711_out0;
assign v$RM_3540_out0 = v$_3063_out0;
assign v$RM_3541_out0 = v$_3873_out0;
assign v$RM_3542_out0 = v$_3835_out0;
assign v$RM_3543_out0 = v$_2167_out0;
assign v$RM_3544_out0 = v$_1785_out0;
assign v$RM_3545_out0 = v$_3151_out0;
assign v$RM_3546_out0 = v$_6812_out0;
assign v$RM_3547_out0 = v$_480_out0;
assign v$RM_3548_out0 = v$_3097_out0;
assign v$RM_3758_out0 = v$_7671_out0;
assign v$RM_3759_out0 = v$_8796_out0;
assign v$RM_3761_out0 = v$_10746_out0;
assign v$RM_3762_out0 = v$_13475_out0;
assign v$RM_3763_out0 = v$_8726_out0;
assign v$RM_3764_out0 = v$_3078_out0;
assign v$RM_3765_out0 = v$_3888_out0;
assign v$RM_3766_out0 = v$_3850_out0;
assign v$RM_3767_out0 = v$_2182_out0;
assign v$RM_3768_out0 = v$_1800_out0;
assign v$RM_3769_out0 = v$_3166_out0;
assign v$RM_3770_out0 = v$_6827_out0;
assign v$RM_3771_out0 = v$_495_out0;
assign v$RM_3772_out0 = v$_3112_out0;
assign v$CIN_9989_out0 = v$_2206_out0;
assign v$CIN_10213_out0 = v$_2220_out0;
assign v$RM_11685_out0 = v$_2514_out0;
assign v$RM_12149_out0 = v$_2529_out0;
assign v$RD_6238_out0 = v$CIN_9989_out0;
assign v$RD_6702_out0 = v$CIN_10213_out0;
assign v$G1_8100_out0 = ((v$RD_6245_out0 && !v$RM_11685_out0) || (!v$RD_6245_out0) && v$RM_11685_out0);
assign v$G1_8564_out0 = ((v$RD_6709_out0 && !v$RM_12149_out0) || (!v$RD_6709_out0) && v$RM_12149_out0);
assign v$RM_11673_out0 = v$RM_3534_out0;
assign v$RM_11675_out0 = v$RM_3535_out0;
assign v$RM_11679_out0 = v$RM_3537_out0;
assign v$RM_11681_out0 = v$RM_3538_out0;
assign v$RM_11683_out0 = v$RM_3539_out0;
assign v$RM_11686_out0 = v$RM_3540_out0;
assign v$RM_11688_out0 = v$RM_3541_out0;
assign v$RM_11690_out0 = v$RM_3542_out0;
assign v$RM_11692_out0 = v$RM_3543_out0;
assign v$RM_11694_out0 = v$RM_3544_out0;
assign v$RM_11696_out0 = v$RM_3545_out0;
assign v$RM_11698_out0 = v$RM_3546_out0;
assign v$RM_11700_out0 = v$RM_3547_out0;
assign v$RM_11702_out0 = v$RM_3548_out0;
assign v$RM_12137_out0 = v$RM_3758_out0;
assign v$RM_12139_out0 = v$RM_3759_out0;
assign v$RM_12143_out0 = v$RM_3761_out0;
assign v$RM_12145_out0 = v$RM_3762_out0;
assign v$RM_12147_out0 = v$RM_3763_out0;
assign v$RM_12150_out0 = v$RM_3764_out0;
assign v$RM_12152_out0 = v$RM_3765_out0;
assign v$RM_12154_out0 = v$RM_3766_out0;
assign v$RM_12156_out0 = v$RM_3767_out0;
assign v$RM_12158_out0 = v$RM_3768_out0;
assign v$RM_12160_out0 = v$RM_3769_out0;
assign v$RM_12162_out0 = v$RM_3770_out0;
assign v$RM_12164_out0 = v$RM_3771_out0;
assign v$RM_12166_out0 = v$RM_3772_out0;
assign v$G2_12636_out0 = v$RD_6245_out0 && v$RM_11685_out0;
assign v$G2_13100_out0 = v$RD_6709_out0 && v$RM_12149_out0;
assign v$CARRY_5245_out0 = v$G2_12636_out0;
assign v$CARRY_5709_out0 = v$G2_13100_out0;
assign v$G1_8088_out0 = ((v$RD_6233_out0 && !v$RM_11673_out0) || (!v$RD_6233_out0) && v$RM_11673_out0);
assign v$G1_8090_out0 = ((v$RD_6235_out0 && !v$RM_11675_out0) || (!v$RD_6235_out0) && v$RM_11675_out0);
assign v$G1_8094_out0 = ((v$RD_6239_out0 && !v$RM_11679_out0) || (!v$RD_6239_out0) && v$RM_11679_out0);
assign v$G1_8096_out0 = ((v$RD_6241_out0 && !v$RM_11681_out0) || (!v$RD_6241_out0) && v$RM_11681_out0);
assign v$G1_8098_out0 = ((v$RD_6243_out0 && !v$RM_11683_out0) || (!v$RD_6243_out0) && v$RM_11683_out0);
assign v$G1_8101_out0 = ((v$RD_6246_out0 && !v$RM_11686_out0) || (!v$RD_6246_out0) && v$RM_11686_out0);
assign v$G1_8103_out0 = ((v$RD_6248_out0 && !v$RM_11688_out0) || (!v$RD_6248_out0) && v$RM_11688_out0);
assign v$G1_8105_out0 = ((v$RD_6250_out0 && !v$RM_11690_out0) || (!v$RD_6250_out0) && v$RM_11690_out0);
assign v$G1_8107_out0 = ((v$RD_6252_out0 && !v$RM_11692_out0) || (!v$RD_6252_out0) && v$RM_11692_out0);
assign v$G1_8109_out0 = ((v$RD_6254_out0 && !v$RM_11694_out0) || (!v$RD_6254_out0) && v$RM_11694_out0);
assign v$G1_8111_out0 = ((v$RD_6256_out0 && !v$RM_11696_out0) || (!v$RD_6256_out0) && v$RM_11696_out0);
assign v$G1_8113_out0 = ((v$RD_6258_out0 && !v$RM_11698_out0) || (!v$RD_6258_out0) && v$RM_11698_out0);
assign v$G1_8115_out0 = ((v$RD_6260_out0 && !v$RM_11700_out0) || (!v$RD_6260_out0) && v$RM_11700_out0);
assign v$G1_8117_out0 = ((v$RD_6262_out0 && !v$RM_11702_out0) || (!v$RD_6262_out0) && v$RM_11702_out0);
assign v$G1_8552_out0 = ((v$RD_6697_out0 && !v$RM_12137_out0) || (!v$RD_6697_out0) && v$RM_12137_out0);
assign v$G1_8554_out0 = ((v$RD_6699_out0 && !v$RM_12139_out0) || (!v$RD_6699_out0) && v$RM_12139_out0);
assign v$G1_8558_out0 = ((v$RD_6703_out0 && !v$RM_12143_out0) || (!v$RD_6703_out0) && v$RM_12143_out0);
assign v$G1_8560_out0 = ((v$RD_6705_out0 && !v$RM_12145_out0) || (!v$RD_6705_out0) && v$RM_12145_out0);
assign v$G1_8562_out0 = ((v$RD_6707_out0 && !v$RM_12147_out0) || (!v$RD_6707_out0) && v$RM_12147_out0);
assign v$G1_8565_out0 = ((v$RD_6710_out0 && !v$RM_12150_out0) || (!v$RD_6710_out0) && v$RM_12150_out0);
assign v$G1_8567_out0 = ((v$RD_6712_out0 && !v$RM_12152_out0) || (!v$RD_6712_out0) && v$RM_12152_out0);
assign v$G1_8569_out0 = ((v$RD_6714_out0 && !v$RM_12154_out0) || (!v$RD_6714_out0) && v$RM_12154_out0);
assign v$G1_8571_out0 = ((v$RD_6716_out0 && !v$RM_12156_out0) || (!v$RD_6716_out0) && v$RM_12156_out0);
assign v$G1_8573_out0 = ((v$RD_6718_out0 && !v$RM_12158_out0) || (!v$RD_6718_out0) && v$RM_12158_out0);
assign v$G1_8575_out0 = ((v$RD_6720_out0 && !v$RM_12160_out0) || (!v$RD_6720_out0) && v$RM_12160_out0);
assign v$G1_8577_out0 = ((v$RD_6722_out0 && !v$RM_12162_out0) || (!v$RD_6722_out0) && v$RM_12162_out0);
assign v$G1_8579_out0 = ((v$RD_6724_out0 && !v$RM_12164_out0) || (!v$RD_6724_out0) && v$RM_12164_out0);
assign v$G1_8581_out0 = ((v$RD_6726_out0 && !v$RM_12166_out0) || (!v$RD_6726_out0) && v$RM_12166_out0);
assign v$S_9246_out0 = v$G1_8100_out0;
assign v$S_9710_out0 = v$G1_8564_out0;
assign v$G2_12624_out0 = v$RD_6233_out0 && v$RM_11673_out0;
assign v$G2_12626_out0 = v$RD_6235_out0 && v$RM_11675_out0;
assign v$G2_12630_out0 = v$RD_6239_out0 && v$RM_11679_out0;
assign v$G2_12632_out0 = v$RD_6241_out0 && v$RM_11681_out0;
assign v$G2_12634_out0 = v$RD_6243_out0 && v$RM_11683_out0;
assign v$G2_12637_out0 = v$RD_6246_out0 && v$RM_11686_out0;
assign v$G2_12639_out0 = v$RD_6248_out0 && v$RM_11688_out0;
assign v$G2_12641_out0 = v$RD_6250_out0 && v$RM_11690_out0;
assign v$G2_12643_out0 = v$RD_6252_out0 && v$RM_11692_out0;
assign v$G2_12645_out0 = v$RD_6254_out0 && v$RM_11694_out0;
assign v$G2_12647_out0 = v$RD_6256_out0 && v$RM_11696_out0;
assign v$G2_12649_out0 = v$RD_6258_out0 && v$RM_11698_out0;
assign v$G2_12651_out0 = v$RD_6260_out0 && v$RM_11700_out0;
assign v$G2_12653_out0 = v$RD_6262_out0 && v$RM_11702_out0;
assign v$G2_13088_out0 = v$RD_6697_out0 && v$RM_12137_out0;
assign v$G2_13090_out0 = v$RD_6699_out0 && v$RM_12139_out0;
assign v$G2_13094_out0 = v$RD_6703_out0 && v$RM_12143_out0;
assign v$G2_13096_out0 = v$RD_6705_out0 && v$RM_12145_out0;
assign v$G2_13098_out0 = v$RD_6707_out0 && v$RM_12147_out0;
assign v$G2_13101_out0 = v$RD_6710_out0 && v$RM_12150_out0;
assign v$G2_13103_out0 = v$RD_6712_out0 && v$RM_12152_out0;
assign v$G2_13105_out0 = v$RD_6714_out0 && v$RM_12154_out0;
assign v$G2_13107_out0 = v$RD_6716_out0 && v$RM_12156_out0;
assign v$G2_13109_out0 = v$RD_6718_out0 && v$RM_12158_out0;
assign v$G2_13111_out0 = v$RD_6720_out0 && v$RM_12160_out0;
assign v$G2_13113_out0 = v$RD_6722_out0 && v$RM_12162_out0;
assign v$G2_13115_out0 = v$RD_6724_out0 && v$RM_12164_out0;
assign v$G2_13117_out0 = v$RD_6726_out0 && v$RM_12166_out0;
assign v$S_4677_out0 = v$S_9246_out0;
assign v$S_4692_out0 = v$S_9710_out0;
assign v$CARRY_5233_out0 = v$G2_12624_out0;
assign v$CARRY_5235_out0 = v$G2_12626_out0;
assign v$CARRY_5239_out0 = v$G2_12630_out0;
assign v$CARRY_5241_out0 = v$G2_12632_out0;
assign v$CARRY_5243_out0 = v$G2_12634_out0;
assign v$CARRY_5246_out0 = v$G2_12637_out0;
assign v$CARRY_5248_out0 = v$G2_12639_out0;
assign v$CARRY_5250_out0 = v$G2_12641_out0;
assign v$CARRY_5252_out0 = v$G2_12643_out0;
assign v$CARRY_5254_out0 = v$G2_12645_out0;
assign v$CARRY_5256_out0 = v$G2_12647_out0;
assign v$CARRY_5258_out0 = v$G2_12649_out0;
assign v$CARRY_5260_out0 = v$G2_12651_out0;
assign v$CARRY_5262_out0 = v$G2_12653_out0;
assign v$CARRY_5697_out0 = v$G2_13088_out0;
assign v$CARRY_5699_out0 = v$G2_13090_out0;
assign v$CARRY_5703_out0 = v$G2_13094_out0;
assign v$CARRY_5705_out0 = v$G2_13096_out0;
assign v$CARRY_5707_out0 = v$G2_13098_out0;
assign v$CARRY_5710_out0 = v$G2_13101_out0;
assign v$CARRY_5712_out0 = v$G2_13103_out0;
assign v$CARRY_5714_out0 = v$G2_13105_out0;
assign v$CARRY_5716_out0 = v$G2_13107_out0;
assign v$CARRY_5718_out0 = v$G2_13109_out0;
assign v$CARRY_5720_out0 = v$G2_13111_out0;
assign v$CARRY_5722_out0 = v$G2_13113_out0;
assign v$CARRY_5724_out0 = v$G2_13115_out0;
assign v$CARRY_5726_out0 = v$G2_13117_out0;
assign v$S_9234_out0 = v$G1_8088_out0;
assign v$S_9236_out0 = v$G1_8090_out0;
assign v$S_9240_out0 = v$G1_8094_out0;
assign v$S_9242_out0 = v$G1_8096_out0;
assign v$S_9244_out0 = v$G1_8098_out0;
assign v$S_9247_out0 = v$G1_8101_out0;
assign v$S_9249_out0 = v$G1_8103_out0;
assign v$S_9251_out0 = v$G1_8105_out0;
assign v$S_9253_out0 = v$G1_8107_out0;
assign v$S_9255_out0 = v$G1_8109_out0;
assign v$S_9257_out0 = v$G1_8111_out0;
assign v$S_9259_out0 = v$G1_8113_out0;
assign v$S_9261_out0 = v$G1_8115_out0;
assign v$S_9263_out0 = v$G1_8117_out0;
assign v$S_9698_out0 = v$G1_8552_out0;
assign v$S_9700_out0 = v$G1_8554_out0;
assign v$S_9704_out0 = v$G1_8558_out0;
assign v$S_9706_out0 = v$G1_8560_out0;
assign v$S_9708_out0 = v$G1_8562_out0;
assign v$S_9711_out0 = v$G1_8565_out0;
assign v$S_9713_out0 = v$G1_8567_out0;
assign v$S_9715_out0 = v$G1_8569_out0;
assign v$S_9717_out0 = v$G1_8571_out0;
assign v$S_9719_out0 = v$G1_8573_out0;
assign v$S_9721_out0 = v$G1_8575_out0;
assign v$S_9723_out0 = v$G1_8577_out0;
assign v$S_9725_out0 = v$G1_8579_out0;
assign v$S_9727_out0 = v$G1_8581_out0;
assign v$CIN_9995_out0 = v$CARRY_5245_out0;
assign v$CIN_10219_out0 = v$CARRY_5709_out0;
assign v$RD_6251_out0 = v$CIN_9995_out0;
assign v$RD_6715_out0 = v$CIN_10219_out0;
assign v$_10767_out0 = { v$_9802_out0,v$S_4677_out0 };
assign v$_10768_out0 = { v$_9803_out0,v$S_4692_out0 };
assign v$RM_11674_out0 = v$S_9234_out0;
assign v$RM_11676_out0 = v$S_9236_out0;
assign v$RM_11680_out0 = v$S_9240_out0;
assign v$RM_11682_out0 = v$S_9242_out0;
assign v$RM_11684_out0 = v$S_9244_out0;
assign v$RM_11687_out0 = v$S_9247_out0;
assign v$RM_11689_out0 = v$S_9249_out0;
assign v$RM_11691_out0 = v$S_9251_out0;
assign v$RM_11693_out0 = v$S_9253_out0;
assign v$RM_11695_out0 = v$S_9255_out0;
assign v$RM_11697_out0 = v$S_9257_out0;
assign v$RM_11699_out0 = v$S_9259_out0;
assign v$RM_11701_out0 = v$S_9261_out0;
assign v$RM_11703_out0 = v$S_9263_out0;
assign v$RM_12138_out0 = v$S_9698_out0;
assign v$RM_12140_out0 = v$S_9700_out0;
assign v$RM_12144_out0 = v$S_9704_out0;
assign v$RM_12146_out0 = v$S_9706_out0;
assign v$RM_12148_out0 = v$S_9708_out0;
assign v$RM_12151_out0 = v$S_9711_out0;
assign v$RM_12153_out0 = v$S_9713_out0;
assign v$RM_12155_out0 = v$S_9715_out0;
assign v$RM_12157_out0 = v$S_9717_out0;
assign v$RM_12159_out0 = v$S_9719_out0;
assign v$RM_12161_out0 = v$S_9721_out0;
assign v$RM_12163_out0 = v$S_9723_out0;
assign v$RM_12165_out0 = v$S_9725_out0;
assign v$RM_12167_out0 = v$S_9727_out0;
assign v$G1_8106_out0 = ((v$RD_6251_out0 && !v$RM_11691_out0) || (!v$RD_6251_out0) && v$RM_11691_out0);
assign v$G1_8570_out0 = ((v$RD_6715_out0 && !v$RM_12155_out0) || (!v$RD_6715_out0) && v$RM_12155_out0);
assign v$G2_12642_out0 = v$RD_6251_out0 && v$RM_11691_out0;
assign v$G2_13106_out0 = v$RD_6715_out0 && v$RM_12155_out0;
assign v$CARRY_5251_out0 = v$G2_12642_out0;
assign v$CARRY_5715_out0 = v$G2_13106_out0;
assign v$S_9252_out0 = v$G1_8106_out0;
assign v$S_9716_out0 = v$G1_8570_out0;
assign v$S_1406_out0 = v$S_9252_out0;
assign v$S_1630_out0 = v$S_9716_out0;
assign v$G1_4182_out0 = v$CARRY_5251_out0 || v$CARRY_5250_out0;
assign v$G1_4406_out0 = v$CARRY_5715_out0 || v$CARRY_5714_out0;
assign v$COUT_874_out0 = v$G1_4182_out0;
assign v$COUT_1098_out0 = v$G1_4406_out0;
assign v$CIN_10001_out0 = v$COUT_874_out0;
assign v$CIN_10225_out0 = v$COUT_1098_out0;
assign v$RD_6263_out0 = v$CIN_10001_out0;
assign v$RD_6727_out0 = v$CIN_10225_out0;
assign v$G1_8118_out0 = ((v$RD_6263_out0 && !v$RM_11703_out0) || (!v$RD_6263_out0) && v$RM_11703_out0);
assign v$G1_8582_out0 = ((v$RD_6727_out0 && !v$RM_12167_out0) || (!v$RD_6727_out0) && v$RM_12167_out0);
assign v$G2_12654_out0 = v$RD_6263_out0 && v$RM_11703_out0;
assign v$G2_13118_out0 = v$RD_6727_out0 && v$RM_12167_out0;
assign v$CARRY_5263_out0 = v$G2_12654_out0;
assign v$CARRY_5727_out0 = v$G2_13118_out0;
assign v$S_9264_out0 = v$G1_8118_out0;
assign v$S_9728_out0 = v$G1_8582_out0;
assign v$S_1412_out0 = v$S_9264_out0;
assign v$S_1636_out0 = v$S_9728_out0;
assign v$G1_4188_out0 = v$CARRY_5263_out0 || v$CARRY_5262_out0;
assign v$G1_4412_out0 = v$CARRY_5727_out0 || v$CARRY_5726_out0;
assign v$COUT_880_out0 = v$G1_4188_out0;
assign v$COUT_1104_out0 = v$G1_4412_out0;
assign v$_4794_out0 = { v$S_1406_out0,v$S_1412_out0 };
assign v$_4809_out0 = { v$S_1630_out0,v$S_1636_out0 };
assign v$CIN_9996_out0 = v$COUT_880_out0;
assign v$CIN_10220_out0 = v$COUT_1104_out0;
assign v$RD_6253_out0 = v$CIN_9996_out0;
assign v$RD_6717_out0 = v$CIN_10220_out0;
assign v$G1_8108_out0 = ((v$RD_6253_out0 && !v$RM_11693_out0) || (!v$RD_6253_out0) && v$RM_11693_out0);
assign v$G1_8572_out0 = ((v$RD_6717_out0 && !v$RM_12157_out0) || (!v$RD_6717_out0) && v$RM_12157_out0);
assign v$G2_12644_out0 = v$RD_6253_out0 && v$RM_11693_out0;
assign v$G2_13108_out0 = v$RD_6717_out0 && v$RM_12157_out0;
assign v$CARRY_5253_out0 = v$G2_12644_out0;
assign v$CARRY_5717_out0 = v$G2_13108_out0;
assign v$S_9254_out0 = v$G1_8108_out0;
assign v$S_9718_out0 = v$G1_8572_out0;
assign v$S_1407_out0 = v$S_9254_out0;
assign v$S_1631_out0 = v$S_9718_out0;
assign v$G1_4183_out0 = v$CARRY_5253_out0 || v$CARRY_5252_out0;
assign v$G1_4407_out0 = v$CARRY_5717_out0 || v$CARRY_5716_out0;
assign v$COUT_875_out0 = v$G1_4183_out0;
assign v$COUT_1099_out0 = v$G1_4407_out0;
assign v$_2564_out0 = { v$_4794_out0,v$S_1407_out0 };
assign v$_2579_out0 = { v$_4809_out0,v$S_1631_out0 };
assign v$CIN_9991_out0 = v$COUT_875_out0;
assign v$CIN_10215_out0 = v$COUT_1099_out0;
assign v$RD_6242_out0 = v$CIN_9991_out0;
assign v$RD_6706_out0 = v$CIN_10215_out0;
assign v$G1_8097_out0 = ((v$RD_6242_out0 && !v$RM_11682_out0) || (!v$RD_6242_out0) && v$RM_11682_out0);
assign v$G1_8561_out0 = ((v$RD_6706_out0 && !v$RM_12146_out0) || (!v$RD_6706_out0) && v$RM_12146_out0);
assign v$G2_12633_out0 = v$RD_6242_out0 && v$RM_11682_out0;
assign v$G2_13097_out0 = v$RD_6706_out0 && v$RM_12146_out0;
assign v$CARRY_5242_out0 = v$G2_12633_out0;
assign v$CARRY_5706_out0 = v$G2_13097_out0;
assign v$S_9243_out0 = v$G1_8097_out0;
assign v$S_9707_out0 = v$G1_8561_out0;
assign v$S_1402_out0 = v$S_9243_out0;
assign v$S_1626_out0 = v$S_9707_out0;
assign v$G1_4178_out0 = v$CARRY_5242_out0 || v$CARRY_5241_out0;
assign v$G1_4402_out0 = v$CARRY_5706_out0 || v$CARRY_5705_out0;
assign v$COUT_870_out0 = v$G1_4178_out0;
assign v$COUT_1094_out0 = v$G1_4402_out0;
assign v$_7044_out0 = { v$_2564_out0,v$S_1402_out0 };
assign v$_7059_out0 = { v$_2579_out0,v$S_1626_out0 };
assign v$CIN_9990_out0 = v$COUT_870_out0;
assign v$CIN_10214_out0 = v$COUT_1094_out0;
assign v$RD_6240_out0 = v$CIN_9990_out0;
assign v$RD_6704_out0 = v$CIN_10214_out0;
assign v$G1_8095_out0 = ((v$RD_6240_out0 && !v$RM_11680_out0) || (!v$RD_6240_out0) && v$RM_11680_out0);
assign v$G1_8559_out0 = ((v$RD_6704_out0 && !v$RM_12144_out0) || (!v$RD_6704_out0) && v$RM_12144_out0);
assign v$G2_12631_out0 = v$RD_6240_out0 && v$RM_11680_out0;
assign v$G2_13095_out0 = v$RD_6704_out0 && v$RM_12144_out0;
assign v$CARRY_5240_out0 = v$G2_12631_out0;
assign v$CARRY_5704_out0 = v$G2_13095_out0;
assign v$S_9241_out0 = v$G1_8095_out0;
assign v$S_9705_out0 = v$G1_8559_out0;
assign v$S_1401_out0 = v$S_9241_out0;
assign v$S_1625_out0 = v$S_9705_out0;
assign v$G1_4177_out0 = v$CARRY_5240_out0 || v$CARRY_5239_out0;
assign v$G1_4401_out0 = v$CARRY_5704_out0 || v$CARRY_5703_out0;
assign v$COUT_869_out0 = v$G1_4177_out0;
assign v$COUT_1093_out0 = v$G1_4401_out0;
assign v$_13530_out0 = { v$_7044_out0,v$S_1401_out0 };
assign v$_13545_out0 = { v$_7059_out0,v$S_1625_out0 };
assign v$CIN_9997_out0 = v$COUT_869_out0;
assign v$CIN_10221_out0 = v$COUT_1093_out0;
assign v$RD_6255_out0 = v$CIN_9997_out0;
assign v$RD_6719_out0 = v$CIN_10221_out0;
assign v$G1_8110_out0 = ((v$RD_6255_out0 && !v$RM_11695_out0) || (!v$RD_6255_out0) && v$RM_11695_out0);
assign v$G1_8574_out0 = ((v$RD_6719_out0 && !v$RM_12159_out0) || (!v$RD_6719_out0) && v$RM_12159_out0);
assign v$G2_12646_out0 = v$RD_6255_out0 && v$RM_11695_out0;
assign v$G2_13110_out0 = v$RD_6719_out0 && v$RM_12159_out0;
assign v$CARRY_5255_out0 = v$G2_12646_out0;
assign v$CARRY_5719_out0 = v$G2_13110_out0;
assign v$S_9256_out0 = v$G1_8110_out0;
assign v$S_9720_out0 = v$G1_8574_out0;
assign v$S_1408_out0 = v$S_9256_out0;
assign v$S_1632_out0 = v$S_9720_out0;
assign v$G1_4184_out0 = v$CARRY_5255_out0 || v$CARRY_5254_out0;
assign v$G1_4408_out0 = v$CARRY_5719_out0 || v$CARRY_5718_out0;
assign v$COUT_876_out0 = v$G1_4184_out0;
assign v$COUT_1100_out0 = v$G1_4408_out0;
assign v$_3323_out0 = { v$_13530_out0,v$S_1408_out0 };
assign v$_3338_out0 = { v$_13545_out0,v$S_1632_out0 };
assign v$CIN_9998_out0 = v$COUT_876_out0;
assign v$CIN_10222_out0 = v$COUT_1100_out0;
assign v$RD_6257_out0 = v$CIN_9998_out0;
assign v$RD_6721_out0 = v$CIN_10222_out0;
assign v$G1_8112_out0 = ((v$RD_6257_out0 && !v$RM_11697_out0) || (!v$RD_6257_out0) && v$RM_11697_out0);
assign v$G1_8576_out0 = ((v$RD_6721_out0 && !v$RM_12161_out0) || (!v$RD_6721_out0) && v$RM_12161_out0);
assign v$G2_12648_out0 = v$RD_6257_out0 && v$RM_11697_out0;
assign v$G2_13112_out0 = v$RD_6721_out0 && v$RM_12161_out0;
assign v$CARRY_5257_out0 = v$G2_12648_out0;
assign v$CARRY_5721_out0 = v$G2_13112_out0;
assign v$S_9258_out0 = v$G1_8112_out0;
assign v$S_9722_out0 = v$G1_8576_out0;
assign v$S_1409_out0 = v$S_9258_out0;
assign v$S_1633_out0 = v$S_9722_out0;
assign v$G1_4185_out0 = v$CARRY_5257_out0 || v$CARRY_5256_out0;
assign v$G1_4409_out0 = v$CARRY_5721_out0 || v$CARRY_5720_out0;
assign v$COUT_877_out0 = v$G1_4185_out0;
assign v$COUT_1101_out0 = v$G1_4409_out0;
assign v$_7159_out0 = { v$_3323_out0,v$S_1409_out0 };
assign v$_7174_out0 = { v$_3338_out0,v$S_1633_out0 };
assign v$CIN_10000_out0 = v$COUT_877_out0;
assign v$CIN_10224_out0 = v$COUT_1101_out0;
assign v$RD_6261_out0 = v$CIN_10000_out0;
assign v$RD_6725_out0 = v$CIN_10224_out0;
assign v$G1_8116_out0 = ((v$RD_6261_out0 && !v$RM_11701_out0) || (!v$RD_6261_out0) && v$RM_11701_out0);
assign v$G1_8580_out0 = ((v$RD_6725_out0 && !v$RM_12165_out0) || (!v$RD_6725_out0) && v$RM_12165_out0);
assign v$G2_12652_out0 = v$RD_6261_out0 && v$RM_11701_out0;
assign v$G2_13116_out0 = v$RD_6725_out0 && v$RM_12165_out0;
assign v$CARRY_5261_out0 = v$G2_12652_out0;
assign v$CARRY_5725_out0 = v$G2_13116_out0;
assign v$S_9262_out0 = v$G1_8116_out0;
assign v$S_9726_out0 = v$G1_8580_out0;
assign v$S_1411_out0 = v$S_9262_out0;
assign v$S_1635_out0 = v$S_9726_out0;
assign v$G1_4187_out0 = v$CARRY_5261_out0 || v$CARRY_5260_out0;
assign v$G1_4411_out0 = v$CARRY_5725_out0 || v$CARRY_5724_out0;
assign v$COUT_879_out0 = v$G1_4187_out0;
assign v$COUT_1103_out0 = v$G1_4411_out0;
assign v$_4761_out0 = { v$_7159_out0,v$S_1411_out0 };
assign v$_4776_out0 = { v$_7174_out0,v$S_1635_out0 };
assign v$CIN_9993_out0 = v$COUT_879_out0;
assign v$CIN_10217_out0 = v$COUT_1103_out0;
assign v$RD_6247_out0 = v$CIN_9993_out0;
assign v$RD_6711_out0 = v$CIN_10217_out0;
assign v$G1_8102_out0 = ((v$RD_6247_out0 && !v$RM_11687_out0) || (!v$RD_6247_out0) && v$RM_11687_out0);
assign v$G1_8566_out0 = ((v$RD_6711_out0 && !v$RM_12151_out0) || (!v$RD_6711_out0) && v$RM_12151_out0);
assign v$G2_12638_out0 = v$RD_6247_out0 && v$RM_11687_out0;
assign v$G2_13102_out0 = v$RD_6711_out0 && v$RM_12151_out0;
assign v$CARRY_5247_out0 = v$G2_12638_out0;
assign v$CARRY_5711_out0 = v$G2_13102_out0;
assign v$S_9248_out0 = v$G1_8102_out0;
assign v$S_9712_out0 = v$G1_8566_out0;
assign v$S_1404_out0 = v$S_9248_out0;
assign v$S_1628_out0 = v$S_9712_out0;
assign v$G1_4180_out0 = v$CARRY_5247_out0 || v$CARRY_5246_out0;
assign v$G1_4404_out0 = v$CARRY_5711_out0 || v$CARRY_5710_out0;
assign v$COUT_872_out0 = v$G1_4180_out0;
assign v$COUT_1096_out0 = v$G1_4404_out0;
assign v$_6938_out0 = { v$_4761_out0,v$S_1404_out0 };
assign v$_6953_out0 = { v$_4776_out0,v$S_1628_out0 };
assign v$CIN_9994_out0 = v$COUT_872_out0;
assign v$CIN_10218_out0 = v$COUT_1096_out0;
assign v$RD_6249_out0 = v$CIN_9994_out0;
assign v$RD_6713_out0 = v$CIN_10218_out0;
assign v$G1_8104_out0 = ((v$RD_6249_out0 && !v$RM_11689_out0) || (!v$RD_6249_out0) && v$RM_11689_out0);
assign v$G1_8568_out0 = ((v$RD_6713_out0 && !v$RM_12153_out0) || (!v$RD_6713_out0) && v$RM_12153_out0);
assign v$G2_12640_out0 = v$RD_6249_out0 && v$RM_11689_out0;
assign v$G2_13104_out0 = v$RD_6713_out0 && v$RM_12153_out0;
assign v$CARRY_5249_out0 = v$G2_12640_out0;
assign v$CARRY_5713_out0 = v$G2_13104_out0;
assign v$S_9250_out0 = v$G1_8104_out0;
assign v$S_9714_out0 = v$G1_8568_out0;
assign v$S_1405_out0 = v$S_9250_out0;
assign v$S_1629_out0 = v$S_9714_out0;
assign v$G1_4181_out0 = v$CARRY_5249_out0 || v$CARRY_5248_out0;
assign v$G1_4405_out0 = v$CARRY_5713_out0 || v$CARRY_5712_out0;
assign v$COUT_873_out0 = v$G1_4181_out0;
assign v$COUT_1097_out0 = v$G1_4405_out0;
assign v$_5814_out0 = { v$_6938_out0,v$S_1405_out0 };
assign v$_5829_out0 = { v$_6953_out0,v$S_1629_out0 };
assign v$CIN_9999_out0 = v$COUT_873_out0;
assign v$CIN_10223_out0 = v$COUT_1097_out0;
assign v$RD_6259_out0 = v$CIN_9999_out0;
assign v$RD_6723_out0 = v$CIN_10223_out0;
assign v$G1_8114_out0 = ((v$RD_6259_out0 && !v$RM_11699_out0) || (!v$RD_6259_out0) && v$RM_11699_out0);
assign v$G1_8578_out0 = ((v$RD_6723_out0 && !v$RM_12163_out0) || (!v$RD_6723_out0) && v$RM_12163_out0);
assign v$G2_12650_out0 = v$RD_6259_out0 && v$RM_11699_out0;
assign v$G2_13114_out0 = v$RD_6723_out0 && v$RM_12163_out0;
assign v$CARRY_5259_out0 = v$G2_12650_out0;
assign v$CARRY_5723_out0 = v$G2_13114_out0;
assign v$S_9260_out0 = v$G1_8114_out0;
assign v$S_9724_out0 = v$G1_8578_out0;
assign v$S_1410_out0 = v$S_9260_out0;
assign v$S_1634_out0 = v$S_9724_out0;
assign v$G1_4186_out0 = v$CARRY_5259_out0 || v$CARRY_5258_out0;
assign v$G1_4410_out0 = v$CARRY_5723_out0 || v$CARRY_5722_out0;
assign v$COUT_878_out0 = v$G1_4186_out0;
assign v$COUT_1102_out0 = v$G1_4410_out0;
assign v$_2038_out0 = { v$_5814_out0,v$S_1410_out0 };
assign v$_2053_out0 = { v$_5829_out0,v$S_1634_out0 };
assign v$CIN_9987_out0 = v$COUT_878_out0;
assign v$CIN_10211_out0 = v$COUT_1102_out0;
assign v$RD_6234_out0 = v$CIN_9987_out0;
assign v$RD_6698_out0 = v$CIN_10211_out0;
assign v$G1_8089_out0 = ((v$RD_6234_out0 && !v$RM_11674_out0) || (!v$RD_6234_out0) && v$RM_11674_out0);
assign v$G1_8553_out0 = ((v$RD_6698_out0 && !v$RM_12138_out0) || (!v$RD_6698_out0) && v$RM_12138_out0);
assign v$G2_12625_out0 = v$RD_6234_out0 && v$RM_11674_out0;
assign v$G2_13089_out0 = v$RD_6698_out0 && v$RM_12138_out0;
assign v$CARRY_5234_out0 = v$G2_12625_out0;
assign v$CARRY_5698_out0 = v$G2_13089_out0;
assign v$S_9235_out0 = v$G1_8089_out0;
assign v$S_9699_out0 = v$G1_8553_out0;
assign v$S_1398_out0 = v$S_9235_out0;
assign v$S_1622_out0 = v$S_9699_out0;
assign v$G1_4174_out0 = v$CARRY_5234_out0 || v$CARRY_5233_out0;
assign v$G1_4398_out0 = v$CARRY_5698_out0 || v$CARRY_5697_out0;
assign v$COUT_866_out0 = v$G1_4174_out0;
assign v$COUT_1090_out0 = v$G1_4398_out0;
assign v$_2805_out0 = { v$_2038_out0,v$S_1398_out0 };
assign v$_2820_out0 = { v$_2053_out0,v$S_1622_out0 };
assign v$CIN_9992_out0 = v$COUT_866_out0;
assign v$CIN_10216_out0 = v$COUT_1090_out0;
assign v$RD_6244_out0 = v$CIN_9992_out0;
assign v$RD_6708_out0 = v$CIN_10216_out0;
assign v$G1_8099_out0 = ((v$RD_6244_out0 && !v$RM_11684_out0) || (!v$RD_6244_out0) && v$RM_11684_out0);
assign v$G1_8563_out0 = ((v$RD_6708_out0 && !v$RM_12148_out0) || (!v$RD_6708_out0) && v$RM_12148_out0);
assign v$G2_12635_out0 = v$RD_6244_out0 && v$RM_11684_out0;
assign v$G2_13099_out0 = v$RD_6708_out0 && v$RM_12148_out0;
assign v$CARRY_5244_out0 = v$G2_12635_out0;
assign v$CARRY_5708_out0 = v$G2_13099_out0;
assign v$S_9245_out0 = v$G1_8099_out0;
assign v$S_9709_out0 = v$G1_8563_out0;
assign v$S_1403_out0 = v$S_9245_out0;
assign v$S_1627_out0 = v$S_9709_out0;
assign v$G1_4179_out0 = v$CARRY_5244_out0 || v$CARRY_5243_out0;
assign v$G1_4403_out0 = v$CARRY_5708_out0 || v$CARRY_5707_out0;
assign v$COUT_871_out0 = v$G1_4179_out0;
assign v$COUT_1095_out0 = v$G1_4403_out0;
assign v$_1837_out0 = { v$_2805_out0,v$S_1403_out0 };
assign v$_1852_out0 = { v$_2820_out0,v$S_1627_out0 };
assign v$CIN_9988_out0 = v$COUT_871_out0;
assign v$CIN_10212_out0 = v$COUT_1095_out0;
assign v$RD_6236_out0 = v$CIN_9988_out0;
assign v$RD_6700_out0 = v$CIN_10212_out0;
assign v$G1_8091_out0 = ((v$RD_6236_out0 && !v$RM_11676_out0) || (!v$RD_6236_out0) && v$RM_11676_out0);
assign v$G1_8555_out0 = ((v$RD_6700_out0 && !v$RM_12140_out0) || (!v$RD_6700_out0) && v$RM_12140_out0);
assign v$G2_12627_out0 = v$RD_6236_out0 && v$RM_11676_out0;
assign v$G2_13091_out0 = v$RD_6700_out0 && v$RM_12140_out0;
assign v$CARRY_5236_out0 = v$G2_12627_out0;
assign v$CARRY_5700_out0 = v$G2_13091_out0;
assign v$S_9237_out0 = v$G1_8091_out0;
assign v$S_9701_out0 = v$G1_8555_out0;
assign v$S_1399_out0 = v$S_9237_out0;
assign v$S_1623_out0 = v$S_9701_out0;
assign v$G1_4175_out0 = v$CARRY_5236_out0 || v$CARRY_5235_out0;
assign v$G1_4399_out0 = v$CARRY_5700_out0 || v$CARRY_5699_out0;
assign v$COUT_867_out0 = v$G1_4175_out0;
assign v$COUT_1091_out0 = v$G1_4399_out0;
assign v$_4561_out0 = { v$_1837_out0,v$S_1399_out0 };
assign v$_4576_out0 = { v$_1852_out0,v$S_1623_out0 };
assign v$RM_3536_out0 = v$COUT_867_out0;
assign v$RM_3760_out0 = v$COUT_1091_out0;
assign v$RM_11677_out0 = v$RM_3536_out0;
assign v$RM_12141_out0 = v$RM_3760_out0;
assign v$G1_8092_out0 = ((v$RD_6237_out0 && !v$RM_11677_out0) || (!v$RD_6237_out0) && v$RM_11677_out0);
assign v$G1_8556_out0 = ((v$RD_6701_out0 && !v$RM_12141_out0) || (!v$RD_6701_out0) && v$RM_12141_out0);
assign v$G2_12628_out0 = v$RD_6237_out0 && v$RM_11677_out0;
assign v$G2_13092_out0 = v$RD_6701_out0 && v$RM_12141_out0;
assign v$CARRY_5237_out0 = v$G2_12628_out0;
assign v$CARRY_5701_out0 = v$G2_13092_out0;
assign v$S_9238_out0 = v$G1_8092_out0;
assign v$S_9702_out0 = v$G1_8556_out0;
assign v$RM_11678_out0 = v$S_9238_out0;
assign v$RM_12142_out0 = v$S_9702_out0;
assign v$G1_8093_out0 = ((v$RD_6238_out0 && !v$RM_11678_out0) || (!v$RD_6238_out0) && v$RM_11678_out0);
assign v$G1_8557_out0 = ((v$RD_6702_out0 && !v$RM_12142_out0) || (!v$RD_6702_out0) && v$RM_12142_out0);
assign v$G2_12629_out0 = v$RD_6238_out0 && v$RM_11678_out0;
assign v$G2_13093_out0 = v$RD_6702_out0 && v$RM_12142_out0;
assign v$CARRY_5238_out0 = v$G2_12629_out0;
assign v$CARRY_5702_out0 = v$G2_13093_out0;
assign v$S_9239_out0 = v$G1_8093_out0;
assign v$S_9703_out0 = v$G1_8557_out0;
assign v$S_1400_out0 = v$S_9239_out0;
assign v$S_1624_out0 = v$S_9703_out0;
assign v$G1_4176_out0 = v$CARRY_5238_out0 || v$CARRY_5237_out0;
assign v$G1_4400_out0 = v$CARRY_5702_out0 || v$CARRY_5701_out0;
assign v$COUT_868_out0 = v$G1_4176_out0;
assign v$COUT_1092_out0 = v$G1_4400_out0;
assign v$_10663_out0 = { v$_4561_out0,v$S_1400_out0 };
assign v$_10678_out0 = { v$_4576_out0,v$S_1624_out0 };
assign v$_10958_out0 = { v$_10663_out0,v$COUT_868_out0 };
assign v$_10973_out0 = { v$_10678_out0,v$COUT_1092_out0 };
assign v$COUT_10928_out0 = v$_10958_out0;
assign v$COUT_10943_out0 = v$_10973_out0;
assign v$CIN_2362_out0 = v$COUT_10928_out0;
assign v$CIN_2377_out0 = v$COUT_10943_out0;
assign v$_475_out0 = v$CIN_2362_out0[8:8];
assign v$_490_out0 = v$CIN_2377_out0[8:8];
assign v$_1780_out0 = v$CIN_2362_out0[6:6];
assign v$_1795_out0 = v$CIN_2377_out0[6:6];
assign v$_2162_out0 = v$CIN_2362_out0[3:3];
assign v$_2177_out0 = v$CIN_2377_out0[3:3];
assign v$_2201_out0 = v$CIN_2362_out0[15:15];
assign v$_2215_out0 = v$CIN_2377_out0[15:15];
assign v$_2509_out0 = v$CIN_2362_out0[0:0];
assign v$_2524_out0 = v$CIN_2377_out0[0:0];
assign v$_3058_out0 = v$CIN_2362_out0[9:9];
assign v$_3073_out0 = v$CIN_2377_out0[9:9];
assign v$_3092_out0 = v$CIN_2362_out0[2:2];
assign v$_3107_out0 = v$CIN_2377_out0[2:2];
assign v$_3146_out0 = v$CIN_2362_out0[7:7];
assign v$_3161_out0 = v$CIN_2377_out0[7:7];
assign v$_3830_out0 = v$CIN_2362_out0[1:1];
assign v$_3845_out0 = v$CIN_2377_out0[1:1];
assign v$_3868_out0 = v$CIN_2362_out0[10:10];
assign v$_3883_out0 = v$CIN_2377_out0[10:10];
assign v$_6807_out0 = v$CIN_2362_out0[11:11];
assign v$_6822_out0 = v$CIN_2377_out0[11:11];
assign v$_7651_out0 = v$CIN_2362_out0[12:12];
assign v$_7666_out0 = v$CIN_2377_out0[12:12];
assign v$_8706_out0 = v$CIN_2362_out0[13:13];
assign v$_8721_out0 = v$CIN_2377_out0[13:13];
assign v$_8776_out0 = v$CIN_2362_out0[14:14];
assign v$_8791_out0 = v$CIN_2377_out0[14:14];
assign v$_10726_out0 = v$CIN_2362_out0[5:5];
assign v$_10741_out0 = v$CIN_2377_out0[5:5];
assign v$_13455_out0 = v$CIN_2362_out0[4:4];
assign v$_13470_out0 = v$CIN_2377_out0[4:4];
assign v$RM_3459_out0 = v$_7651_out0;
assign v$RM_3460_out0 = v$_8776_out0;
assign v$RM_3462_out0 = v$_10726_out0;
assign v$RM_3463_out0 = v$_13455_out0;
assign v$RM_3464_out0 = v$_8706_out0;
assign v$RM_3465_out0 = v$_3058_out0;
assign v$RM_3466_out0 = v$_3868_out0;
assign v$RM_3467_out0 = v$_3830_out0;
assign v$RM_3468_out0 = v$_2162_out0;
assign v$RM_3469_out0 = v$_1780_out0;
assign v$RM_3470_out0 = v$_3146_out0;
assign v$RM_3471_out0 = v$_6807_out0;
assign v$RM_3472_out0 = v$_475_out0;
assign v$RM_3473_out0 = v$_3092_out0;
assign v$RM_3683_out0 = v$_7666_out0;
assign v$RM_3684_out0 = v$_8791_out0;
assign v$RM_3686_out0 = v$_10741_out0;
assign v$RM_3687_out0 = v$_13470_out0;
assign v$RM_3688_out0 = v$_8721_out0;
assign v$RM_3689_out0 = v$_3073_out0;
assign v$RM_3690_out0 = v$_3883_out0;
assign v$RM_3691_out0 = v$_3845_out0;
assign v$RM_3692_out0 = v$_2177_out0;
assign v$RM_3693_out0 = v$_1795_out0;
assign v$RM_3694_out0 = v$_3161_out0;
assign v$RM_3695_out0 = v$_6822_out0;
assign v$RM_3696_out0 = v$_490_out0;
assign v$RM_3697_out0 = v$_3107_out0;
assign v$CIN_9914_out0 = v$_2201_out0;
assign v$CIN_10138_out0 = v$_2215_out0;
assign v$RM_11530_out0 = v$_2509_out0;
assign v$RM_11994_out0 = v$_2524_out0;
assign v$RD_6083_out0 = v$CIN_9914_out0;
assign v$RD_6547_out0 = v$CIN_10138_out0;
assign v$G1_7945_out0 = ((v$RD_6090_out0 && !v$RM_11530_out0) || (!v$RD_6090_out0) && v$RM_11530_out0);
assign v$G1_8409_out0 = ((v$RD_6554_out0 && !v$RM_11994_out0) || (!v$RD_6554_out0) && v$RM_11994_out0);
assign v$RM_11518_out0 = v$RM_3459_out0;
assign v$RM_11520_out0 = v$RM_3460_out0;
assign v$RM_11524_out0 = v$RM_3462_out0;
assign v$RM_11526_out0 = v$RM_3463_out0;
assign v$RM_11528_out0 = v$RM_3464_out0;
assign v$RM_11531_out0 = v$RM_3465_out0;
assign v$RM_11533_out0 = v$RM_3466_out0;
assign v$RM_11535_out0 = v$RM_3467_out0;
assign v$RM_11537_out0 = v$RM_3468_out0;
assign v$RM_11539_out0 = v$RM_3469_out0;
assign v$RM_11541_out0 = v$RM_3470_out0;
assign v$RM_11543_out0 = v$RM_3471_out0;
assign v$RM_11545_out0 = v$RM_3472_out0;
assign v$RM_11547_out0 = v$RM_3473_out0;
assign v$RM_11982_out0 = v$RM_3683_out0;
assign v$RM_11984_out0 = v$RM_3684_out0;
assign v$RM_11988_out0 = v$RM_3686_out0;
assign v$RM_11990_out0 = v$RM_3687_out0;
assign v$RM_11992_out0 = v$RM_3688_out0;
assign v$RM_11995_out0 = v$RM_3689_out0;
assign v$RM_11997_out0 = v$RM_3690_out0;
assign v$RM_11999_out0 = v$RM_3691_out0;
assign v$RM_12001_out0 = v$RM_3692_out0;
assign v$RM_12003_out0 = v$RM_3693_out0;
assign v$RM_12005_out0 = v$RM_3694_out0;
assign v$RM_12007_out0 = v$RM_3695_out0;
assign v$RM_12009_out0 = v$RM_3696_out0;
assign v$RM_12011_out0 = v$RM_3697_out0;
assign v$G2_12481_out0 = v$RD_6090_out0 && v$RM_11530_out0;
assign v$G2_12945_out0 = v$RD_6554_out0 && v$RM_11994_out0;
assign v$CARRY_5090_out0 = v$G2_12481_out0;
assign v$CARRY_5554_out0 = v$G2_12945_out0;
assign v$G1_7933_out0 = ((v$RD_6078_out0 && !v$RM_11518_out0) || (!v$RD_6078_out0) && v$RM_11518_out0);
assign v$G1_7935_out0 = ((v$RD_6080_out0 && !v$RM_11520_out0) || (!v$RD_6080_out0) && v$RM_11520_out0);
assign v$G1_7939_out0 = ((v$RD_6084_out0 && !v$RM_11524_out0) || (!v$RD_6084_out0) && v$RM_11524_out0);
assign v$G1_7941_out0 = ((v$RD_6086_out0 && !v$RM_11526_out0) || (!v$RD_6086_out0) && v$RM_11526_out0);
assign v$G1_7943_out0 = ((v$RD_6088_out0 && !v$RM_11528_out0) || (!v$RD_6088_out0) && v$RM_11528_out0);
assign v$G1_7946_out0 = ((v$RD_6091_out0 && !v$RM_11531_out0) || (!v$RD_6091_out0) && v$RM_11531_out0);
assign v$G1_7948_out0 = ((v$RD_6093_out0 && !v$RM_11533_out0) || (!v$RD_6093_out0) && v$RM_11533_out0);
assign v$G1_7950_out0 = ((v$RD_6095_out0 && !v$RM_11535_out0) || (!v$RD_6095_out0) && v$RM_11535_out0);
assign v$G1_7952_out0 = ((v$RD_6097_out0 && !v$RM_11537_out0) || (!v$RD_6097_out0) && v$RM_11537_out0);
assign v$G1_7954_out0 = ((v$RD_6099_out0 && !v$RM_11539_out0) || (!v$RD_6099_out0) && v$RM_11539_out0);
assign v$G1_7956_out0 = ((v$RD_6101_out0 && !v$RM_11541_out0) || (!v$RD_6101_out0) && v$RM_11541_out0);
assign v$G1_7958_out0 = ((v$RD_6103_out0 && !v$RM_11543_out0) || (!v$RD_6103_out0) && v$RM_11543_out0);
assign v$G1_7960_out0 = ((v$RD_6105_out0 && !v$RM_11545_out0) || (!v$RD_6105_out0) && v$RM_11545_out0);
assign v$G1_7962_out0 = ((v$RD_6107_out0 && !v$RM_11547_out0) || (!v$RD_6107_out0) && v$RM_11547_out0);
assign v$G1_8397_out0 = ((v$RD_6542_out0 && !v$RM_11982_out0) || (!v$RD_6542_out0) && v$RM_11982_out0);
assign v$G1_8399_out0 = ((v$RD_6544_out0 && !v$RM_11984_out0) || (!v$RD_6544_out0) && v$RM_11984_out0);
assign v$G1_8403_out0 = ((v$RD_6548_out0 && !v$RM_11988_out0) || (!v$RD_6548_out0) && v$RM_11988_out0);
assign v$G1_8405_out0 = ((v$RD_6550_out0 && !v$RM_11990_out0) || (!v$RD_6550_out0) && v$RM_11990_out0);
assign v$G1_8407_out0 = ((v$RD_6552_out0 && !v$RM_11992_out0) || (!v$RD_6552_out0) && v$RM_11992_out0);
assign v$G1_8410_out0 = ((v$RD_6555_out0 && !v$RM_11995_out0) || (!v$RD_6555_out0) && v$RM_11995_out0);
assign v$G1_8412_out0 = ((v$RD_6557_out0 && !v$RM_11997_out0) || (!v$RD_6557_out0) && v$RM_11997_out0);
assign v$G1_8414_out0 = ((v$RD_6559_out0 && !v$RM_11999_out0) || (!v$RD_6559_out0) && v$RM_11999_out0);
assign v$G1_8416_out0 = ((v$RD_6561_out0 && !v$RM_12001_out0) || (!v$RD_6561_out0) && v$RM_12001_out0);
assign v$G1_8418_out0 = ((v$RD_6563_out0 && !v$RM_12003_out0) || (!v$RD_6563_out0) && v$RM_12003_out0);
assign v$G1_8420_out0 = ((v$RD_6565_out0 && !v$RM_12005_out0) || (!v$RD_6565_out0) && v$RM_12005_out0);
assign v$G1_8422_out0 = ((v$RD_6567_out0 && !v$RM_12007_out0) || (!v$RD_6567_out0) && v$RM_12007_out0);
assign v$G1_8424_out0 = ((v$RD_6569_out0 && !v$RM_12009_out0) || (!v$RD_6569_out0) && v$RM_12009_out0);
assign v$G1_8426_out0 = ((v$RD_6571_out0 && !v$RM_12011_out0) || (!v$RD_6571_out0) && v$RM_12011_out0);
assign v$S_9091_out0 = v$G1_7945_out0;
assign v$S_9555_out0 = v$G1_8409_out0;
assign v$G2_12469_out0 = v$RD_6078_out0 && v$RM_11518_out0;
assign v$G2_12471_out0 = v$RD_6080_out0 && v$RM_11520_out0;
assign v$G2_12475_out0 = v$RD_6084_out0 && v$RM_11524_out0;
assign v$G2_12477_out0 = v$RD_6086_out0 && v$RM_11526_out0;
assign v$G2_12479_out0 = v$RD_6088_out0 && v$RM_11528_out0;
assign v$G2_12482_out0 = v$RD_6091_out0 && v$RM_11531_out0;
assign v$G2_12484_out0 = v$RD_6093_out0 && v$RM_11533_out0;
assign v$G2_12486_out0 = v$RD_6095_out0 && v$RM_11535_out0;
assign v$G2_12488_out0 = v$RD_6097_out0 && v$RM_11537_out0;
assign v$G2_12490_out0 = v$RD_6099_out0 && v$RM_11539_out0;
assign v$G2_12492_out0 = v$RD_6101_out0 && v$RM_11541_out0;
assign v$G2_12494_out0 = v$RD_6103_out0 && v$RM_11543_out0;
assign v$G2_12496_out0 = v$RD_6105_out0 && v$RM_11545_out0;
assign v$G2_12498_out0 = v$RD_6107_out0 && v$RM_11547_out0;
assign v$G2_12933_out0 = v$RD_6542_out0 && v$RM_11982_out0;
assign v$G2_12935_out0 = v$RD_6544_out0 && v$RM_11984_out0;
assign v$G2_12939_out0 = v$RD_6548_out0 && v$RM_11988_out0;
assign v$G2_12941_out0 = v$RD_6550_out0 && v$RM_11990_out0;
assign v$G2_12943_out0 = v$RD_6552_out0 && v$RM_11992_out0;
assign v$G2_12946_out0 = v$RD_6555_out0 && v$RM_11995_out0;
assign v$G2_12948_out0 = v$RD_6557_out0 && v$RM_11997_out0;
assign v$G2_12950_out0 = v$RD_6559_out0 && v$RM_11999_out0;
assign v$G2_12952_out0 = v$RD_6561_out0 && v$RM_12001_out0;
assign v$G2_12954_out0 = v$RD_6563_out0 && v$RM_12003_out0;
assign v$G2_12956_out0 = v$RD_6565_out0 && v$RM_12005_out0;
assign v$G2_12958_out0 = v$RD_6567_out0 && v$RM_12007_out0;
assign v$G2_12960_out0 = v$RD_6569_out0 && v$RM_12009_out0;
assign v$G2_12962_out0 = v$RD_6571_out0 && v$RM_12011_out0;
assign v$S_4672_out0 = v$S_9091_out0;
assign v$S_4687_out0 = v$S_9555_out0;
assign v$CARRY_5078_out0 = v$G2_12469_out0;
assign v$CARRY_5080_out0 = v$G2_12471_out0;
assign v$CARRY_5084_out0 = v$G2_12475_out0;
assign v$CARRY_5086_out0 = v$G2_12477_out0;
assign v$CARRY_5088_out0 = v$G2_12479_out0;
assign v$CARRY_5091_out0 = v$G2_12482_out0;
assign v$CARRY_5093_out0 = v$G2_12484_out0;
assign v$CARRY_5095_out0 = v$G2_12486_out0;
assign v$CARRY_5097_out0 = v$G2_12488_out0;
assign v$CARRY_5099_out0 = v$G2_12490_out0;
assign v$CARRY_5101_out0 = v$G2_12492_out0;
assign v$CARRY_5103_out0 = v$G2_12494_out0;
assign v$CARRY_5105_out0 = v$G2_12496_out0;
assign v$CARRY_5107_out0 = v$G2_12498_out0;
assign v$CARRY_5542_out0 = v$G2_12933_out0;
assign v$CARRY_5544_out0 = v$G2_12935_out0;
assign v$CARRY_5548_out0 = v$G2_12939_out0;
assign v$CARRY_5550_out0 = v$G2_12941_out0;
assign v$CARRY_5552_out0 = v$G2_12943_out0;
assign v$CARRY_5555_out0 = v$G2_12946_out0;
assign v$CARRY_5557_out0 = v$G2_12948_out0;
assign v$CARRY_5559_out0 = v$G2_12950_out0;
assign v$CARRY_5561_out0 = v$G2_12952_out0;
assign v$CARRY_5563_out0 = v$G2_12954_out0;
assign v$CARRY_5565_out0 = v$G2_12956_out0;
assign v$CARRY_5567_out0 = v$G2_12958_out0;
assign v$CARRY_5569_out0 = v$G2_12960_out0;
assign v$CARRY_5571_out0 = v$G2_12962_out0;
assign v$S_9079_out0 = v$G1_7933_out0;
assign v$S_9081_out0 = v$G1_7935_out0;
assign v$S_9085_out0 = v$G1_7939_out0;
assign v$S_9087_out0 = v$G1_7941_out0;
assign v$S_9089_out0 = v$G1_7943_out0;
assign v$S_9092_out0 = v$G1_7946_out0;
assign v$S_9094_out0 = v$G1_7948_out0;
assign v$S_9096_out0 = v$G1_7950_out0;
assign v$S_9098_out0 = v$G1_7952_out0;
assign v$S_9100_out0 = v$G1_7954_out0;
assign v$S_9102_out0 = v$G1_7956_out0;
assign v$S_9104_out0 = v$G1_7958_out0;
assign v$S_9106_out0 = v$G1_7960_out0;
assign v$S_9108_out0 = v$G1_7962_out0;
assign v$S_9543_out0 = v$G1_8397_out0;
assign v$S_9545_out0 = v$G1_8399_out0;
assign v$S_9549_out0 = v$G1_8403_out0;
assign v$S_9551_out0 = v$G1_8405_out0;
assign v$S_9553_out0 = v$G1_8407_out0;
assign v$S_9556_out0 = v$G1_8410_out0;
assign v$S_9558_out0 = v$G1_8412_out0;
assign v$S_9560_out0 = v$G1_8414_out0;
assign v$S_9562_out0 = v$G1_8416_out0;
assign v$S_9564_out0 = v$G1_8418_out0;
assign v$S_9566_out0 = v$G1_8420_out0;
assign v$S_9568_out0 = v$G1_8422_out0;
assign v$S_9570_out0 = v$G1_8424_out0;
assign v$S_9572_out0 = v$G1_8426_out0;
assign v$CIN_9920_out0 = v$CARRY_5090_out0;
assign v$CIN_10144_out0 = v$CARRY_5554_out0;
assign v$RD_6096_out0 = v$CIN_9920_out0;
assign v$RD_6560_out0 = v$CIN_10144_out0;
assign v$RM_11519_out0 = v$S_9079_out0;
assign v$RM_11521_out0 = v$S_9081_out0;
assign v$RM_11525_out0 = v$S_9085_out0;
assign v$RM_11527_out0 = v$S_9087_out0;
assign v$RM_11529_out0 = v$S_9089_out0;
assign v$RM_11532_out0 = v$S_9092_out0;
assign v$RM_11534_out0 = v$S_9094_out0;
assign v$RM_11536_out0 = v$S_9096_out0;
assign v$RM_11538_out0 = v$S_9098_out0;
assign v$RM_11540_out0 = v$S_9100_out0;
assign v$RM_11542_out0 = v$S_9102_out0;
assign v$RM_11544_out0 = v$S_9104_out0;
assign v$RM_11546_out0 = v$S_9106_out0;
assign v$RM_11548_out0 = v$S_9108_out0;
assign v$RM_11983_out0 = v$S_9543_out0;
assign v$RM_11985_out0 = v$S_9545_out0;
assign v$RM_11989_out0 = v$S_9549_out0;
assign v$RM_11991_out0 = v$S_9551_out0;
assign v$RM_11993_out0 = v$S_9553_out0;
assign v$RM_11996_out0 = v$S_9556_out0;
assign v$RM_11998_out0 = v$S_9558_out0;
assign v$RM_12000_out0 = v$S_9560_out0;
assign v$RM_12002_out0 = v$S_9562_out0;
assign v$RM_12004_out0 = v$S_9564_out0;
assign v$RM_12006_out0 = v$S_9566_out0;
assign v$RM_12008_out0 = v$S_9568_out0;
assign v$RM_12010_out0 = v$S_9570_out0;
assign v$RM_12012_out0 = v$S_9572_out0;
assign v$_13709_out0 = { v$_10767_out0,v$S_4672_out0 };
assign v$_13710_out0 = { v$_10768_out0,v$S_4687_out0 };
assign v$G1_7951_out0 = ((v$RD_6096_out0 && !v$RM_11536_out0) || (!v$RD_6096_out0) && v$RM_11536_out0);
assign v$G1_8415_out0 = ((v$RD_6560_out0 && !v$RM_12000_out0) || (!v$RD_6560_out0) && v$RM_12000_out0);
assign v$G2_12487_out0 = v$RD_6096_out0 && v$RM_11536_out0;
assign v$G2_12951_out0 = v$RD_6560_out0 && v$RM_12000_out0;
assign v$CARRY_5096_out0 = v$G2_12487_out0;
assign v$CARRY_5560_out0 = v$G2_12951_out0;
assign v$S_9097_out0 = v$G1_7951_out0;
assign v$S_9561_out0 = v$G1_8415_out0;
assign v$S_1331_out0 = v$S_9097_out0;
assign v$S_1555_out0 = v$S_9561_out0;
assign v$G1_4107_out0 = v$CARRY_5096_out0 || v$CARRY_5095_out0;
assign v$G1_4331_out0 = v$CARRY_5560_out0 || v$CARRY_5559_out0;
assign v$COUT_799_out0 = v$G1_4107_out0;
assign v$COUT_1023_out0 = v$G1_4331_out0;
assign v$CIN_9926_out0 = v$COUT_799_out0;
assign v$CIN_10150_out0 = v$COUT_1023_out0;
assign v$RD_6108_out0 = v$CIN_9926_out0;
assign v$RD_6572_out0 = v$CIN_10150_out0;
assign v$G1_7963_out0 = ((v$RD_6108_out0 && !v$RM_11548_out0) || (!v$RD_6108_out0) && v$RM_11548_out0);
assign v$G1_8427_out0 = ((v$RD_6572_out0 && !v$RM_12012_out0) || (!v$RD_6572_out0) && v$RM_12012_out0);
assign v$G2_12499_out0 = v$RD_6108_out0 && v$RM_11548_out0;
assign v$G2_12963_out0 = v$RD_6572_out0 && v$RM_12012_out0;
assign v$CARRY_5108_out0 = v$G2_12499_out0;
assign v$CARRY_5572_out0 = v$G2_12963_out0;
assign v$S_9109_out0 = v$G1_7963_out0;
assign v$S_9573_out0 = v$G1_8427_out0;
assign v$S_1337_out0 = v$S_9109_out0;
assign v$S_1561_out0 = v$S_9573_out0;
assign v$G1_4113_out0 = v$CARRY_5108_out0 || v$CARRY_5107_out0;
assign v$G1_4337_out0 = v$CARRY_5572_out0 || v$CARRY_5571_out0;
assign v$COUT_805_out0 = v$G1_4113_out0;
assign v$COUT_1029_out0 = v$G1_4337_out0;
assign v$_4789_out0 = { v$S_1331_out0,v$S_1337_out0 };
assign v$_4804_out0 = { v$S_1555_out0,v$S_1561_out0 };
assign v$CIN_9921_out0 = v$COUT_805_out0;
assign v$CIN_10145_out0 = v$COUT_1029_out0;
assign v$RD_6098_out0 = v$CIN_9921_out0;
assign v$RD_6562_out0 = v$CIN_10145_out0;
assign v$G1_7953_out0 = ((v$RD_6098_out0 && !v$RM_11538_out0) || (!v$RD_6098_out0) && v$RM_11538_out0);
assign v$G1_8417_out0 = ((v$RD_6562_out0 && !v$RM_12002_out0) || (!v$RD_6562_out0) && v$RM_12002_out0);
assign v$G2_12489_out0 = v$RD_6098_out0 && v$RM_11538_out0;
assign v$G2_12953_out0 = v$RD_6562_out0 && v$RM_12002_out0;
assign v$CARRY_5098_out0 = v$G2_12489_out0;
assign v$CARRY_5562_out0 = v$G2_12953_out0;
assign v$S_9099_out0 = v$G1_7953_out0;
assign v$S_9563_out0 = v$G1_8417_out0;
assign v$S_1332_out0 = v$S_9099_out0;
assign v$S_1556_out0 = v$S_9563_out0;
assign v$G1_4108_out0 = v$CARRY_5098_out0 || v$CARRY_5097_out0;
assign v$G1_4332_out0 = v$CARRY_5562_out0 || v$CARRY_5561_out0;
assign v$COUT_800_out0 = v$G1_4108_out0;
assign v$COUT_1024_out0 = v$G1_4332_out0;
assign v$_2559_out0 = { v$_4789_out0,v$S_1332_out0 };
assign v$_2574_out0 = { v$_4804_out0,v$S_1556_out0 };
assign v$CIN_9916_out0 = v$COUT_800_out0;
assign v$CIN_10140_out0 = v$COUT_1024_out0;
assign v$RD_6087_out0 = v$CIN_9916_out0;
assign v$RD_6551_out0 = v$CIN_10140_out0;
assign v$G1_7942_out0 = ((v$RD_6087_out0 && !v$RM_11527_out0) || (!v$RD_6087_out0) && v$RM_11527_out0);
assign v$G1_8406_out0 = ((v$RD_6551_out0 && !v$RM_11991_out0) || (!v$RD_6551_out0) && v$RM_11991_out0);
assign v$G2_12478_out0 = v$RD_6087_out0 && v$RM_11527_out0;
assign v$G2_12942_out0 = v$RD_6551_out0 && v$RM_11991_out0;
assign v$CARRY_5087_out0 = v$G2_12478_out0;
assign v$CARRY_5551_out0 = v$G2_12942_out0;
assign v$S_9088_out0 = v$G1_7942_out0;
assign v$S_9552_out0 = v$G1_8406_out0;
assign v$S_1327_out0 = v$S_9088_out0;
assign v$S_1551_out0 = v$S_9552_out0;
assign v$G1_4103_out0 = v$CARRY_5087_out0 || v$CARRY_5086_out0;
assign v$G1_4327_out0 = v$CARRY_5551_out0 || v$CARRY_5550_out0;
assign v$COUT_795_out0 = v$G1_4103_out0;
assign v$COUT_1019_out0 = v$G1_4327_out0;
assign v$_7039_out0 = { v$_2559_out0,v$S_1327_out0 };
assign v$_7054_out0 = { v$_2574_out0,v$S_1551_out0 };
assign v$CIN_9915_out0 = v$COUT_795_out0;
assign v$CIN_10139_out0 = v$COUT_1019_out0;
assign v$RD_6085_out0 = v$CIN_9915_out0;
assign v$RD_6549_out0 = v$CIN_10139_out0;
assign v$G1_7940_out0 = ((v$RD_6085_out0 && !v$RM_11525_out0) || (!v$RD_6085_out0) && v$RM_11525_out0);
assign v$G1_8404_out0 = ((v$RD_6549_out0 && !v$RM_11989_out0) || (!v$RD_6549_out0) && v$RM_11989_out0);
assign v$G2_12476_out0 = v$RD_6085_out0 && v$RM_11525_out0;
assign v$G2_12940_out0 = v$RD_6549_out0 && v$RM_11989_out0;
assign v$CARRY_5085_out0 = v$G2_12476_out0;
assign v$CARRY_5549_out0 = v$G2_12940_out0;
assign v$S_9086_out0 = v$G1_7940_out0;
assign v$S_9550_out0 = v$G1_8404_out0;
assign v$S_1326_out0 = v$S_9086_out0;
assign v$S_1550_out0 = v$S_9550_out0;
assign v$G1_4102_out0 = v$CARRY_5085_out0 || v$CARRY_5084_out0;
assign v$G1_4326_out0 = v$CARRY_5549_out0 || v$CARRY_5548_out0;
assign v$COUT_794_out0 = v$G1_4102_out0;
assign v$COUT_1018_out0 = v$G1_4326_out0;
assign v$_13525_out0 = { v$_7039_out0,v$S_1326_out0 };
assign v$_13540_out0 = { v$_7054_out0,v$S_1550_out0 };
assign v$CIN_9922_out0 = v$COUT_794_out0;
assign v$CIN_10146_out0 = v$COUT_1018_out0;
assign v$RD_6100_out0 = v$CIN_9922_out0;
assign v$RD_6564_out0 = v$CIN_10146_out0;
assign v$G1_7955_out0 = ((v$RD_6100_out0 && !v$RM_11540_out0) || (!v$RD_6100_out0) && v$RM_11540_out0);
assign v$G1_8419_out0 = ((v$RD_6564_out0 && !v$RM_12004_out0) || (!v$RD_6564_out0) && v$RM_12004_out0);
assign v$G2_12491_out0 = v$RD_6100_out0 && v$RM_11540_out0;
assign v$G2_12955_out0 = v$RD_6564_out0 && v$RM_12004_out0;
assign v$CARRY_5100_out0 = v$G2_12491_out0;
assign v$CARRY_5564_out0 = v$G2_12955_out0;
assign v$S_9101_out0 = v$G1_7955_out0;
assign v$S_9565_out0 = v$G1_8419_out0;
assign v$S_1333_out0 = v$S_9101_out0;
assign v$S_1557_out0 = v$S_9565_out0;
assign v$G1_4109_out0 = v$CARRY_5100_out0 || v$CARRY_5099_out0;
assign v$G1_4333_out0 = v$CARRY_5564_out0 || v$CARRY_5563_out0;
assign v$COUT_801_out0 = v$G1_4109_out0;
assign v$COUT_1025_out0 = v$G1_4333_out0;
assign v$_3318_out0 = { v$_13525_out0,v$S_1333_out0 };
assign v$_3333_out0 = { v$_13540_out0,v$S_1557_out0 };
assign v$CIN_9923_out0 = v$COUT_801_out0;
assign v$CIN_10147_out0 = v$COUT_1025_out0;
assign v$RD_6102_out0 = v$CIN_9923_out0;
assign v$RD_6566_out0 = v$CIN_10147_out0;
assign v$G1_7957_out0 = ((v$RD_6102_out0 && !v$RM_11542_out0) || (!v$RD_6102_out0) && v$RM_11542_out0);
assign v$G1_8421_out0 = ((v$RD_6566_out0 && !v$RM_12006_out0) || (!v$RD_6566_out0) && v$RM_12006_out0);
assign v$G2_12493_out0 = v$RD_6102_out0 && v$RM_11542_out0;
assign v$G2_12957_out0 = v$RD_6566_out0 && v$RM_12006_out0;
assign v$CARRY_5102_out0 = v$G2_12493_out0;
assign v$CARRY_5566_out0 = v$G2_12957_out0;
assign v$S_9103_out0 = v$G1_7957_out0;
assign v$S_9567_out0 = v$G1_8421_out0;
assign v$S_1334_out0 = v$S_9103_out0;
assign v$S_1558_out0 = v$S_9567_out0;
assign v$G1_4110_out0 = v$CARRY_5102_out0 || v$CARRY_5101_out0;
assign v$G1_4334_out0 = v$CARRY_5566_out0 || v$CARRY_5565_out0;
assign v$COUT_802_out0 = v$G1_4110_out0;
assign v$COUT_1026_out0 = v$G1_4334_out0;
assign v$_7154_out0 = { v$_3318_out0,v$S_1334_out0 };
assign v$_7169_out0 = { v$_3333_out0,v$S_1558_out0 };
assign v$CIN_9925_out0 = v$COUT_802_out0;
assign v$CIN_10149_out0 = v$COUT_1026_out0;
assign v$RD_6106_out0 = v$CIN_9925_out0;
assign v$RD_6570_out0 = v$CIN_10149_out0;
assign v$G1_7961_out0 = ((v$RD_6106_out0 && !v$RM_11546_out0) || (!v$RD_6106_out0) && v$RM_11546_out0);
assign v$G1_8425_out0 = ((v$RD_6570_out0 && !v$RM_12010_out0) || (!v$RD_6570_out0) && v$RM_12010_out0);
assign v$G2_12497_out0 = v$RD_6106_out0 && v$RM_11546_out0;
assign v$G2_12961_out0 = v$RD_6570_out0 && v$RM_12010_out0;
assign v$CARRY_5106_out0 = v$G2_12497_out0;
assign v$CARRY_5570_out0 = v$G2_12961_out0;
assign v$S_9107_out0 = v$G1_7961_out0;
assign v$S_9571_out0 = v$G1_8425_out0;
assign v$S_1336_out0 = v$S_9107_out0;
assign v$S_1560_out0 = v$S_9571_out0;
assign v$G1_4112_out0 = v$CARRY_5106_out0 || v$CARRY_5105_out0;
assign v$G1_4336_out0 = v$CARRY_5570_out0 || v$CARRY_5569_out0;
assign v$COUT_804_out0 = v$G1_4112_out0;
assign v$COUT_1028_out0 = v$G1_4336_out0;
assign v$_4756_out0 = { v$_7154_out0,v$S_1336_out0 };
assign v$_4771_out0 = { v$_7169_out0,v$S_1560_out0 };
assign v$CIN_9918_out0 = v$COUT_804_out0;
assign v$CIN_10142_out0 = v$COUT_1028_out0;
assign v$RD_6092_out0 = v$CIN_9918_out0;
assign v$RD_6556_out0 = v$CIN_10142_out0;
assign v$G1_7947_out0 = ((v$RD_6092_out0 && !v$RM_11532_out0) || (!v$RD_6092_out0) && v$RM_11532_out0);
assign v$G1_8411_out0 = ((v$RD_6556_out0 && !v$RM_11996_out0) || (!v$RD_6556_out0) && v$RM_11996_out0);
assign v$G2_12483_out0 = v$RD_6092_out0 && v$RM_11532_out0;
assign v$G2_12947_out0 = v$RD_6556_out0 && v$RM_11996_out0;
assign v$CARRY_5092_out0 = v$G2_12483_out0;
assign v$CARRY_5556_out0 = v$G2_12947_out0;
assign v$S_9093_out0 = v$G1_7947_out0;
assign v$S_9557_out0 = v$G1_8411_out0;
assign v$S_1329_out0 = v$S_9093_out0;
assign v$S_1553_out0 = v$S_9557_out0;
assign v$G1_4105_out0 = v$CARRY_5092_out0 || v$CARRY_5091_out0;
assign v$G1_4329_out0 = v$CARRY_5556_out0 || v$CARRY_5555_out0;
assign v$COUT_797_out0 = v$G1_4105_out0;
assign v$COUT_1021_out0 = v$G1_4329_out0;
assign v$_6933_out0 = { v$_4756_out0,v$S_1329_out0 };
assign v$_6948_out0 = { v$_4771_out0,v$S_1553_out0 };
assign v$CIN_9919_out0 = v$COUT_797_out0;
assign v$CIN_10143_out0 = v$COUT_1021_out0;
assign v$RD_6094_out0 = v$CIN_9919_out0;
assign v$RD_6558_out0 = v$CIN_10143_out0;
assign v$G1_7949_out0 = ((v$RD_6094_out0 && !v$RM_11534_out0) || (!v$RD_6094_out0) && v$RM_11534_out0);
assign v$G1_8413_out0 = ((v$RD_6558_out0 && !v$RM_11998_out0) || (!v$RD_6558_out0) && v$RM_11998_out0);
assign v$G2_12485_out0 = v$RD_6094_out0 && v$RM_11534_out0;
assign v$G2_12949_out0 = v$RD_6558_out0 && v$RM_11998_out0;
assign v$CARRY_5094_out0 = v$G2_12485_out0;
assign v$CARRY_5558_out0 = v$G2_12949_out0;
assign v$S_9095_out0 = v$G1_7949_out0;
assign v$S_9559_out0 = v$G1_8413_out0;
assign v$S_1330_out0 = v$S_9095_out0;
assign v$S_1554_out0 = v$S_9559_out0;
assign v$G1_4106_out0 = v$CARRY_5094_out0 || v$CARRY_5093_out0;
assign v$G1_4330_out0 = v$CARRY_5558_out0 || v$CARRY_5557_out0;
assign v$COUT_798_out0 = v$G1_4106_out0;
assign v$COUT_1022_out0 = v$G1_4330_out0;
assign v$_5809_out0 = { v$_6933_out0,v$S_1330_out0 };
assign v$_5824_out0 = { v$_6948_out0,v$S_1554_out0 };
assign v$CIN_9924_out0 = v$COUT_798_out0;
assign v$CIN_10148_out0 = v$COUT_1022_out0;
assign v$RD_6104_out0 = v$CIN_9924_out0;
assign v$RD_6568_out0 = v$CIN_10148_out0;
assign v$G1_7959_out0 = ((v$RD_6104_out0 && !v$RM_11544_out0) || (!v$RD_6104_out0) && v$RM_11544_out0);
assign v$G1_8423_out0 = ((v$RD_6568_out0 && !v$RM_12008_out0) || (!v$RD_6568_out0) && v$RM_12008_out0);
assign v$G2_12495_out0 = v$RD_6104_out0 && v$RM_11544_out0;
assign v$G2_12959_out0 = v$RD_6568_out0 && v$RM_12008_out0;
assign v$CARRY_5104_out0 = v$G2_12495_out0;
assign v$CARRY_5568_out0 = v$G2_12959_out0;
assign v$S_9105_out0 = v$G1_7959_out0;
assign v$S_9569_out0 = v$G1_8423_out0;
assign v$S_1335_out0 = v$S_9105_out0;
assign v$S_1559_out0 = v$S_9569_out0;
assign v$G1_4111_out0 = v$CARRY_5104_out0 || v$CARRY_5103_out0;
assign v$G1_4335_out0 = v$CARRY_5568_out0 || v$CARRY_5567_out0;
assign v$COUT_803_out0 = v$G1_4111_out0;
assign v$COUT_1027_out0 = v$G1_4335_out0;
assign v$_2033_out0 = { v$_5809_out0,v$S_1335_out0 };
assign v$_2048_out0 = { v$_5824_out0,v$S_1559_out0 };
assign v$CIN_9912_out0 = v$COUT_803_out0;
assign v$CIN_10136_out0 = v$COUT_1027_out0;
assign v$RD_6079_out0 = v$CIN_9912_out0;
assign v$RD_6543_out0 = v$CIN_10136_out0;
assign v$G1_7934_out0 = ((v$RD_6079_out0 && !v$RM_11519_out0) || (!v$RD_6079_out0) && v$RM_11519_out0);
assign v$G1_8398_out0 = ((v$RD_6543_out0 && !v$RM_11983_out0) || (!v$RD_6543_out0) && v$RM_11983_out0);
assign v$G2_12470_out0 = v$RD_6079_out0 && v$RM_11519_out0;
assign v$G2_12934_out0 = v$RD_6543_out0 && v$RM_11983_out0;
assign v$CARRY_5079_out0 = v$G2_12470_out0;
assign v$CARRY_5543_out0 = v$G2_12934_out0;
assign v$S_9080_out0 = v$G1_7934_out0;
assign v$S_9544_out0 = v$G1_8398_out0;
assign v$S_1323_out0 = v$S_9080_out0;
assign v$S_1547_out0 = v$S_9544_out0;
assign v$G1_4099_out0 = v$CARRY_5079_out0 || v$CARRY_5078_out0;
assign v$G1_4323_out0 = v$CARRY_5543_out0 || v$CARRY_5542_out0;
assign v$COUT_791_out0 = v$G1_4099_out0;
assign v$COUT_1015_out0 = v$G1_4323_out0;
assign v$_2800_out0 = { v$_2033_out0,v$S_1323_out0 };
assign v$_2815_out0 = { v$_2048_out0,v$S_1547_out0 };
assign v$CIN_9917_out0 = v$COUT_791_out0;
assign v$CIN_10141_out0 = v$COUT_1015_out0;
assign v$RD_6089_out0 = v$CIN_9917_out0;
assign v$RD_6553_out0 = v$CIN_10141_out0;
assign v$G1_7944_out0 = ((v$RD_6089_out0 && !v$RM_11529_out0) || (!v$RD_6089_out0) && v$RM_11529_out0);
assign v$G1_8408_out0 = ((v$RD_6553_out0 && !v$RM_11993_out0) || (!v$RD_6553_out0) && v$RM_11993_out0);
assign v$G2_12480_out0 = v$RD_6089_out0 && v$RM_11529_out0;
assign v$G2_12944_out0 = v$RD_6553_out0 && v$RM_11993_out0;
assign v$CARRY_5089_out0 = v$G2_12480_out0;
assign v$CARRY_5553_out0 = v$G2_12944_out0;
assign v$S_9090_out0 = v$G1_7944_out0;
assign v$S_9554_out0 = v$G1_8408_out0;
assign v$S_1328_out0 = v$S_9090_out0;
assign v$S_1552_out0 = v$S_9554_out0;
assign v$G1_4104_out0 = v$CARRY_5089_out0 || v$CARRY_5088_out0;
assign v$G1_4328_out0 = v$CARRY_5553_out0 || v$CARRY_5552_out0;
assign v$COUT_796_out0 = v$G1_4104_out0;
assign v$COUT_1020_out0 = v$G1_4328_out0;
assign v$_1832_out0 = { v$_2800_out0,v$S_1328_out0 };
assign v$_1847_out0 = { v$_2815_out0,v$S_1552_out0 };
assign v$CIN_9913_out0 = v$COUT_796_out0;
assign v$CIN_10137_out0 = v$COUT_1020_out0;
assign v$RD_6081_out0 = v$CIN_9913_out0;
assign v$RD_6545_out0 = v$CIN_10137_out0;
assign v$G1_7936_out0 = ((v$RD_6081_out0 && !v$RM_11521_out0) || (!v$RD_6081_out0) && v$RM_11521_out0);
assign v$G1_8400_out0 = ((v$RD_6545_out0 && !v$RM_11985_out0) || (!v$RD_6545_out0) && v$RM_11985_out0);
assign v$G2_12472_out0 = v$RD_6081_out0 && v$RM_11521_out0;
assign v$G2_12936_out0 = v$RD_6545_out0 && v$RM_11985_out0;
assign v$CARRY_5081_out0 = v$G2_12472_out0;
assign v$CARRY_5545_out0 = v$G2_12936_out0;
assign v$S_9082_out0 = v$G1_7936_out0;
assign v$S_9546_out0 = v$G1_8400_out0;
assign v$S_1324_out0 = v$S_9082_out0;
assign v$S_1548_out0 = v$S_9546_out0;
assign v$G1_4100_out0 = v$CARRY_5081_out0 || v$CARRY_5080_out0;
assign v$G1_4324_out0 = v$CARRY_5545_out0 || v$CARRY_5544_out0;
assign v$COUT_792_out0 = v$G1_4100_out0;
assign v$COUT_1016_out0 = v$G1_4324_out0;
assign v$_4556_out0 = { v$_1832_out0,v$S_1324_out0 };
assign v$_4571_out0 = { v$_1847_out0,v$S_1548_out0 };
assign v$RM_3461_out0 = v$COUT_792_out0;
assign v$RM_3685_out0 = v$COUT_1016_out0;
assign v$RM_11522_out0 = v$RM_3461_out0;
assign v$RM_11986_out0 = v$RM_3685_out0;
assign v$G1_7937_out0 = ((v$RD_6082_out0 && !v$RM_11522_out0) || (!v$RD_6082_out0) && v$RM_11522_out0);
assign v$G1_8401_out0 = ((v$RD_6546_out0 && !v$RM_11986_out0) || (!v$RD_6546_out0) && v$RM_11986_out0);
assign v$G2_12473_out0 = v$RD_6082_out0 && v$RM_11522_out0;
assign v$G2_12937_out0 = v$RD_6546_out0 && v$RM_11986_out0;
assign v$CARRY_5082_out0 = v$G2_12473_out0;
assign v$CARRY_5546_out0 = v$G2_12937_out0;
assign v$S_9083_out0 = v$G1_7937_out0;
assign v$S_9547_out0 = v$G1_8401_out0;
assign v$RM_11523_out0 = v$S_9083_out0;
assign v$RM_11987_out0 = v$S_9547_out0;
assign v$G1_7938_out0 = ((v$RD_6083_out0 && !v$RM_11523_out0) || (!v$RD_6083_out0) && v$RM_11523_out0);
assign v$G1_8402_out0 = ((v$RD_6547_out0 && !v$RM_11987_out0) || (!v$RD_6547_out0) && v$RM_11987_out0);
assign v$G2_12474_out0 = v$RD_6083_out0 && v$RM_11523_out0;
assign v$G2_12938_out0 = v$RD_6547_out0 && v$RM_11987_out0;
assign v$CARRY_5083_out0 = v$G2_12474_out0;
assign v$CARRY_5547_out0 = v$G2_12938_out0;
assign v$S_9084_out0 = v$G1_7938_out0;
assign v$S_9548_out0 = v$G1_8402_out0;
assign v$S_1325_out0 = v$S_9084_out0;
assign v$S_1549_out0 = v$S_9548_out0;
assign v$G1_4101_out0 = v$CARRY_5083_out0 || v$CARRY_5082_out0;
assign v$G1_4325_out0 = v$CARRY_5547_out0 || v$CARRY_5546_out0;
assign v$COUT_793_out0 = v$G1_4101_out0;
assign v$COUT_1017_out0 = v$G1_4325_out0;
assign v$_10658_out0 = { v$_4556_out0,v$S_1325_out0 };
assign v$_10673_out0 = { v$_4571_out0,v$S_1549_out0 };
assign v$_10953_out0 = { v$_10658_out0,v$COUT_793_out0 };
assign v$_10968_out0 = { v$_10673_out0,v$COUT_1017_out0 };
assign v$COUT_10923_out0 = v$_10953_out0;
assign v$COUT_10938_out0 = v$_10968_out0;
assign v$CIN_2361_out0 = v$COUT_10923_out0;
assign v$CIN_2376_out0 = v$COUT_10938_out0;
assign v$_474_out0 = v$CIN_2361_out0[8:8];
assign v$_489_out0 = v$CIN_2376_out0[8:8];
assign v$_1779_out0 = v$CIN_2361_out0[6:6];
assign v$_1794_out0 = v$CIN_2376_out0[6:6];
assign v$_2161_out0 = v$CIN_2361_out0[3:3];
assign v$_2176_out0 = v$CIN_2376_out0[3:3];
assign v$_2200_out0 = v$CIN_2361_out0[15:15];
assign v$_2214_out0 = v$CIN_2376_out0[15:15];
assign v$_2508_out0 = v$CIN_2361_out0[0:0];
assign v$_2523_out0 = v$CIN_2376_out0[0:0];
assign v$_3057_out0 = v$CIN_2361_out0[9:9];
assign v$_3072_out0 = v$CIN_2376_out0[9:9];
assign v$_3091_out0 = v$CIN_2361_out0[2:2];
assign v$_3106_out0 = v$CIN_2376_out0[2:2];
assign v$_3145_out0 = v$CIN_2361_out0[7:7];
assign v$_3160_out0 = v$CIN_2376_out0[7:7];
assign v$_3829_out0 = v$CIN_2361_out0[1:1];
assign v$_3844_out0 = v$CIN_2376_out0[1:1];
assign v$_3867_out0 = v$CIN_2361_out0[10:10];
assign v$_3882_out0 = v$CIN_2376_out0[10:10];
assign v$_6806_out0 = v$CIN_2361_out0[11:11];
assign v$_6821_out0 = v$CIN_2376_out0[11:11];
assign v$_7650_out0 = v$CIN_2361_out0[12:12];
assign v$_7665_out0 = v$CIN_2376_out0[12:12];
assign v$_8705_out0 = v$CIN_2361_out0[13:13];
assign v$_8720_out0 = v$CIN_2376_out0[13:13];
assign v$_8775_out0 = v$CIN_2361_out0[14:14];
assign v$_8790_out0 = v$CIN_2376_out0[14:14];
assign v$_10725_out0 = v$CIN_2361_out0[5:5];
assign v$_10740_out0 = v$CIN_2376_out0[5:5];
assign v$_13454_out0 = v$CIN_2361_out0[4:4];
assign v$_13469_out0 = v$CIN_2376_out0[4:4];
assign v$RM_3444_out0 = v$_7650_out0;
assign v$RM_3445_out0 = v$_8775_out0;
assign v$RM_3447_out0 = v$_10725_out0;
assign v$RM_3448_out0 = v$_13454_out0;
assign v$RM_3449_out0 = v$_8705_out0;
assign v$RM_3450_out0 = v$_3057_out0;
assign v$RM_3451_out0 = v$_3867_out0;
assign v$RM_3452_out0 = v$_3829_out0;
assign v$RM_3453_out0 = v$_2161_out0;
assign v$RM_3454_out0 = v$_1779_out0;
assign v$RM_3455_out0 = v$_3145_out0;
assign v$RM_3456_out0 = v$_6806_out0;
assign v$RM_3457_out0 = v$_474_out0;
assign v$RM_3458_out0 = v$_3091_out0;
assign v$RM_3668_out0 = v$_7665_out0;
assign v$RM_3669_out0 = v$_8790_out0;
assign v$RM_3671_out0 = v$_10740_out0;
assign v$RM_3672_out0 = v$_13469_out0;
assign v$RM_3673_out0 = v$_8720_out0;
assign v$RM_3674_out0 = v$_3072_out0;
assign v$RM_3675_out0 = v$_3882_out0;
assign v$RM_3676_out0 = v$_3844_out0;
assign v$RM_3677_out0 = v$_2176_out0;
assign v$RM_3678_out0 = v$_1794_out0;
assign v$RM_3679_out0 = v$_3160_out0;
assign v$RM_3680_out0 = v$_6821_out0;
assign v$RM_3681_out0 = v$_489_out0;
assign v$RM_3682_out0 = v$_3106_out0;
assign v$CIN_9899_out0 = v$_2200_out0;
assign v$CIN_10123_out0 = v$_2214_out0;
assign v$RM_11499_out0 = v$_2508_out0;
assign v$RM_11963_out0 = v$_2523_out0;
assign v$RD_6052_out0 = v$CIN_9899_out0;
assign v$RD_6516_out0 = v$CIN_10123_out0;
assign v$G1_7914_out0 = ((v$RD_6059_out0 && !v$RM_11499_out0) || (!v$RD_6059_out0) && v$RM_11499_out0);
assign v$G1_8378_out0 = ((v$RD_6523_out0 && !v$RM_11963_out0) || (!v$RD_6523_out0) && v$RM_11963_out0);
assign v$RM_11487_out0 = v$RM_3444_out0;
assign v$RM_11489_out0 = v$RM_3445_out0;
assign v$RM_11493_out0 = v$RM_3447_out0;
assign v$RM_11495_out0 = v$RM_3448_out0;
assign v$RM_11497_out0 = v$RM_3449_out0;
assign v$RM_11500_out0 = v$RM_3450_out0;
assign v$RM_11502_out0 = v$RM_3451_out0;
assign v$RM_11504_out0 = v$RM_3452_out0;
assign v$RM_11506_out0 = v$RM_3453_out0;
assign v$RM_11508_out0 = v$RM_3454_out0;
assign v$RM_11510_out0 = v$RM_3455_out0;
assign v$RM_11512_out0 = v$RM_3456_out0;
assign v$RM_11514_out0 = v$RM_3457_out0;
assign v$RM_11516_out0 = v$RM_3458_out0;
assign v$RM_11951_out0 = v$RM_3668_out0;
assign v$RM_11953_out0 = v$RM_3669_out0;
assign v$RM_11957_out0 = v$RM_3671_out0;
assign v$RM_11959_out0 = v$RM_3672_out0;
assign v$RM_11961_out0 = v$RM_3673_out0;
assign v$RM_11964_out0 = v$RM_3674_out0;
assign v$RM_11966_out0 = v$RM_3675_out0;
assign v$RM_11968_out0 = v$RM_3676_out0;
assign v$RM_11970_out0 = v$RM_3677_out0;
assign v$RM_11972_out0 = v$RM_3678_out0;
assign v$RM_11974_out0 = v$RM_3679_out0;
assign v$RM_11976_out0 = v$RM_3680_out0;
assign v$RM_11978_out0 = v$RM_3681_out0;
assign v$RM_11980_out0 = v$RM_3682_out0;
assign v$G2_12450_out0 = v$RD_6059_out0 && v$RM_11499_out0;
assign v$G2_12914_out0 = v$RD_6523_out0 && v$RM_11963_out0;
assign v$CARRY_5059_out0 = v$G2_12450_out0;
assign v$CARRY_5523_out0 = v$G2_12914_out0;
assign v$G1_7902_out0 = ((v$RD_6047_out0 && !v$RM_11487_out0) || (!v$RD_6047_out0) && v$RM_11487_out0);
assign v$G1_7904_out0 = ((v$RD_6049_out0 && !v$RM_11489_out0) || (!v$RD_6049_out0) && v$RM_11489_out0);
assign v$G1_7908_out0 = ((v$RD_6053_out0 && !v$RM_11493_out0) || (!v$RD_6053_out0) && v$RM_11493_out0);
assign v$G1_7910_out0 = ((v$RD_6055_out0 && !v$RM_11495_out0) || (!v$RD_6055_out0) && v$RM_11495_out0);
assign v$G1_7912_out0 = ((v$RD_6057_out0 && !v$RM_11497_out0) || (!v$RD_6057_out0) && v$RM_11497_out0);
assign v$G1_7915_out0 = ((v$RD_6060_out0 && !v$RM_11500_out0) || (!v$RD_6060_out0) && v$RM_11500_out0);
assign v$G1_7917_out0 = ((v$RD_6062_out0 && !v$RM_11502_out0) || (!v$RD_6062_out0) && v$RM_11502_out0);
assign v$G1_7919_out0 = ((v$RD_6064_out0 && !v$RM_11504_out0) || (!v$RD_6064_out0) && v$RM_11504_out0);
assign v$G1_7921_out0 = ((v$RD_6066_out0 && !v$RM_11506_out0) || (!v$RD_6066_out0) && v$RM_11506_out0);
assign v$G1_7923_out0 = ((v$RD_6068_out0 && !v$RM_11508_out0) || (!v$RD_6068_out0) && v$RM_11508_out0);
assign v$G1_7925_out0 = ((v$RD_6070_out0 && !v$RM_11510_out0) || (!v$RD_6070_out0) && v$RM_11510_out0);
assign v$G1_7927_out0 = ((v$RD_6072_out0 && !v$RM_11512_out0) || (!v$RD_6072_out0) && v$RM_11512_out0);
assign v$G1_7929_out0 = ((v$RD_6074_out0 && !v$RM_11514_out0) || (!v$RD_6074_out0) && v$RM_11514_out0);
assign v$G1_7931_out0 = ((v$RD_6076_out0 && !v$RM_11516_out0) || (!v$RD_6076_out0) && v$RM_11516_out0);
assign v$G1_8366_out0 = ((v$RD_6511_out0 && !v$RM_11951_out0) || (!v$RD_6511_out0) && v$RM_11951_out0);
assign v$G1_8368_out0 = ((v$RD_6513_out0 && !v$RM_11953_out0) || (!v$RD_6513_out0) && v$RM_11953_out0);
assign v$G1_8372_out0 = ((v$RD_6517_out0 && !v$RM_11957_out0) || (!v$RD_6517_out0) && v$RM_11957_out0);
assign v$G1_8374_out0 = ((v$RD_6519_out0 && !v$RM_11959_out0) || (!v$RD_6519_out0) && v$RM_11959_out0);
assign v$G1_8376_out0 = ((v$RD_6521_out0 && !v$RM_11961_out0) || (!v$RD_6521_out0) && v$RM_11961_out0);
assign v$G1_8379_out0 = ((v$RD_6524_out0 && !v$RM_11964_out0) || (!v$RD_6524_out0) && v$RM_11964_out0);
assign v$G1_8381_out0 = ((v$RD_6526_out0 && !v$RM_11966_out0) || (!v$RD_6526_out0) && v$RM_11966_out0);
assign v$G1_8383_out0 = ((v$RD_6528_out0 && !v$RM_11968_out0) || (!v$RD_6528_out0) && v$RM_11968_out0);
assign v$G1_8385_out0 = ((v$RD_6530_out0 && !v$RM_11970_out0) || (!v$RD_6530_out0) && v$RM_11970_out0);
assign v$G1_8387_out0 = ((v$RD_6532_out0 && !v$RM_11972_out0) || (!v$RD_6532_out0) && v$RM_11972_out0);
assign v$G1_8389_out0 = ((v$RD_6534_out0 && !v$RM_11974_out0) || (!v$RD_6534_out0) && v$RM_11974_out0);
assign v$G1_8391_out0 = ((v$RD_6536_out0 && !v$RM_11976_out0) || (!v$RD_6536_out0) && v$RM_11976_out0);
assign v$G1_8393_out0 = ((v$RD_6538_out0 && !v$RM_11978_out0) || (!v$RD_6538_out0) && v$RM_11978_out0);
assign v$G1_8395_out0 = ((v$RD_6540_out0 && !v$RM_11980_out0) || (!v$RD_6540_out0) && v$RM_11980_out0);
assign v$S_9060_out0 = v$G1_7914_out0;
assign v$S_9524_out0 = v$G1_8378_out0;
assign v$G2_12438_out0 = v$RD_6047_out0 && v$RM_11487_out0;
assign v$G2_12440_out0 = v$RD_6049_out0 && v$RM_11489_out0;
assign v$G2_12444_out0 = v$RD_6053_out0 && v$RM_11493_out0;
assign v$G2_12446_out0 = v$RD_6055_out0 && v$RM_11495_out0;
assign v$G2_12448_out0 = v$RD_6057_out0 && v$RM_11497_out0;
assign v$G2_12451_out0 = v$RD_6060_out0 && v$RM_11500_out0;
assign v$G2_12453_out0 = v$RD_6062_out0 && v$RM_11502_out0;
assign v$G2_12455_out0 = v$RD_6064_out0 && v$RM_11504_out0;
assign v$G2_12457_out0 = v$RD_6066_out0 && v$RM_11506_out0;
assign v$G2_12459_out0 = v$RD_6068_out0 && v$RM_11508_out0;
assign v$G2_12461_out0 = v$RD_6070_out0 && v$RM_11510_out0;
assign v$G2_12463_out0 = v$RD_6072_out0 && v$RM_11512_out0;
assign v$G2_12465_out0 = v$RD_6074_out0 && v$RM_11514_out0;
assign v$G2_12467_out0 = v$RD_6076_out0 && v$RM_11516_out0;
assign v$G2_12902_out0 = v$RD_6511_out0 && v$RM_11951_out0;
assign v$G2_12904_out0 = v$RD_6513_out0 && v$RM_11953_out0;
assign v$G2_12908_out0 = v$RD_6517_out0 && v$RM_11957_out0;
assign v$G2_12910_out0 = v$RD_6519_out0 && v$RM_11959_out0;
assign v$G2_12912_out0 = v$RD_6521_out0 && v$RM_11961_out0;
assign v$G2_12915_out0 = v$RD_6524_out0 && v$RM_11964_out0;
assign v$G2_12917_out0 = v$RD_6526_out0 && v$RM_11966_out0;
assign v$G2_12919_out0 = v$RD_6528_out0 && v$RM_11968_out0;
assign v$G2_12921_out0 = v$RD_6530_out0 && v$RM_11970_out0;
assign v$G2_12923_out0 = v$RD_6532_out0 && v$RM_11972_out0;
assign v$G2_12925_out0 = v$RD_6534_out0 && v$RM_11974_out0;
assign v$G2_12927_out0 = v$RD_6536_out0 && v$RM_11976_out0;
assign v$G2_12929_out0 = v$RD_6538_out0 && v$RM_11978_out0;
assign v$G2_12931_out0 = v$RD_6540_out0 && v$RM_11980_out0;
assign v$S_4671_out0 = v$S_9060_out0;
assign v$S_4686_out0 = v$S_9524_out0;
assign v$CARRY_5047_out0 = v$G2_12438_out0;
assign v$CARRY_5049_out0 = v$G2_12440_out0;
assign v$CARRY_5053_out0 = v$G2_12444_out0;
assign v$CARRY_5055_out0 = v$G2_12446_out0;
assign v$CARRY_5057_out0 = v$G2_12448_out0;
assign v$CARRY_5060_out0 = v$G2_12451_out0;
assign v$CARRY_5062_out0 = v$G2_12453_out0;
assign v$CARRY_5064_out0 = v$G2_12455_out0;
assign v$CARRY_5066_out0 = v$G2_12457_out0;
assign v$CARRY_5068_out0 = v$G2_12459_out0;
assign v$CARRY_5070_out0 = v$G2_12461_out0;
assign v$CARRY_5072_out0 = v$G2_12463_out0;
assign v$CARRY_5074_out0 = v$G2_12465_out0;
assign v$CARRY_5076_out0 = v$G2_12467_out0;
assign v$CARRY_5511_out0 = v$G2_12902_out0;
assign v$CARRY_5513_out0 = v$G2_12904_out0;
assign v$CARRY_5517_out0 = v$G2_12908_out0;
assign v$CARRY_5519_out0 = v$G2_12910_out0;
assign v$CARRY_5521_out0 = v$G2_12912_out0;
assign v$CARRY_5524_out0 = v$G2_12915_out0;
assign v$CARRY_5526_out0 = v$G2_12917_out0;
assign v$CARRY_5528_out0 = v$G2_12919_out0;
assign v$CARRY_5530_out0 = v$G2_12921_out0;
assign v$CARRY_5532_out0 = v$G2_12923_out0;
assign v$CARRY_5534_out0 = v$G2_12925_out0;
assign v$CARRY_5536_out0 = v$G2_12927_out0;
assign v$CARRY_5538_out0 = v$G2_12929_out0;
assign v$CARRY_5540_out0 = v$G2_12931_out0;
assign v$S_9048_out0 = v$G1_7902_out0;
assign v$S_9050_out0 = v$G1_7904_out0;
assign v$S_9054_out0 = v$G1_7908_out0;
assign v$S_9056_out0 = v$G1_7910_out0;
assign v$S_9058_out0 = v$G1_7912_out0;
assign v$S_9061_out0 = v$G1_7915_out0;
assign v$S_9063_out0 = v$G1_7917_out0;
assign v$S_9065_out0 = v$G1_7919_out0;
assign v$S_9067_out0 = v$G1_7921_out0;
assign v$S_9069_out0 = v$G1_7923_out0;
assign v$S_9071_out0 = v$G1_7925_out0;
assign v$S_9073_out0 = v$G1_7927_out0;
assign v$S_9075_out0 = v$G1_7929_out0;
assign v$S_9077_out0 = v$G1_7931_out0;
assign v$S_9512_out0 = v$G1_8366_out0;
assign v$S_9514_out0 = v$G1_8368_out0;
assign v$S_9518_out0 = v$G1_8372_out0;
assign v$S_9520_out0 = v$G1_8374_out0;
assign v$S_9522_out0 = v$G1_8376_out0;
assign v$S_9525_out0 = v$G1_8379_out0;
assign v$S_9527_out0 = v$G1_8381_out0;
assign v$S_9529_out0 = v$G1_8383_out0;
assign v$S_9531_out0 = v$G1_8385_out0;
assign v$S_9533_out0 = v$G1_8387_out0;
assign v$S_9535_out0 = v$G1_8389_out0;
assign v$S_9537_out0 = v$G1_8391_out0;
assign v$S_9539_out0 = v$G1_8393_out0;
assign v$S_9541_out0 = v$G1_8395_out0;
assign v$CIN_9905_out0 = v$CARRY_5059_out0;
assign v$CIN_10129_out0 = v$CARRY_5523_out0;
assign v$_403_out0 = { v$_13709_out0,v$S_4671_out0 };
assign v$_404_out0 = { v$_13710_out0,v$S_4686_out0 };
assign v$RD_6065_out0 = v$CIN_9905_out0;
assign v$RD_6529_out0 = v$CIN_10129_out0;
assign v$RM_11488_out0 = v$S_9048_out0;
assign v$RM_11490_out0 = v$S_9050_out0;
assign v$RM_11494_out0 = v$S_9054_out0;
assign v$RM_11496_out0 = v$S_9056_out0;
assign v$RM_11498_out0 = v$S_9058_out0;
assign v$RM_11501_out0 = v$S_9061_out0;
assign v$RM_11503_out0 = v$S_9063_out0;
assign v$RM_11505_out0 = v$S_9065_out0;
assign v$RM_11507_out0 = v$S_9067_out0;
assign v$RM_11509_out0 = v$S_9069_out0;
assign v$RM_11511_out0 = v$S_9071_out0;
assign v$RM_11513_out0 = v$S_9073_out0;
assign v$RM_11515_out0 = v$S_9075_out0;
assign v$RM_11517_out0 = v$S_9077_out0;
assign v$RM_11952_out0 = v$S_9512_out0;
assign v$RM_11954_out0 = v$S_9514_out0;
assign v$RM_11958_out0 = v$S_9518_out0;
assign v$RM_11960_out0 = v$S_9520_out0;
assign v$RM_11962_out0 = v$S_9522_out0;
assign v$RM_11965_out0 = v$S_9525_out0;
assign v$RM_11967_out0 = v$S_9527_out0;
assign v$RM_11969_out0 = v$S_9529_out0;
assign v$RM_11971_out0 = v$S_9531_out0;
assign v$RM_11973_out0 = v$S_9533_out0;
assign v$RM_11975_out0 = v$S_9535_out0;
assign v$RM_11977_out0 = v$S_9537_out0;
assign v$RM_11979_out0 = v$S_9539_out0;
assign v$RM_11981_out0 = v$S_9541_out0;
assign v$MUX1_2717_out0 = v$EXEC2_3241_out0 ? v$REG1_13338_out0 : v$_403_out0;
assign v$MUX1_2718_out0 = v$EXEC2_3242_out0 ? v$REG1_13339_out0 : v$_404_out0;
assign v$G1_7920_out0 = ((v$RD_6065_out0 && !v$RM_11505_out0) || (!v$RD_6065_out0) && v$RM_11505_out0);
assign v$G1_8384_out0 = ((v$RD_6529_out0 && !v$RM_11969_out0) || (!v$RD_6529_out0) && v$RM_11969_out0);
assign v$G2_12456_out0 = v$RD_6065_out0 && v$RM_11505_out0;
assign v$G2_12920_out0 = v$RD_6529_out0 && v$RM_11969_out0;
assign v$M$REGIN_271_out0 = v$MUX1_2717_out0;
assign v$M$REGIN_272_out0 = v$MUX1_2718_out0;
assign v$CARRY_5065_out0 = v$G2_12456_out0;
assign v$CARRY_5529_out0 = v$G2_12920_out0;
assign v$S_9066_out0 = v$G1_7920_out0;
assign v$S_9530_out0 = v$G1_8384_out0;
assign v$S_1316_out0 = v$S_9066_out0;
assign v$S_1540_out0 = v$S_9530_out0;
assign v$MULTI$REGIN_2870_out0 = v$M$REGIN_271_out0;
assign v$MULTI$REGIN_2871_out0 = v$M$REGIN_272_out0;
assign v$G1_4092_out0 = v$CARRY_5065_out0 || v$CARRY_5064_out0;
assign v$G1_4316_out0 = v$CARRY_5529_out0 || v$CARRY_5528_out0;
assign v$COUT_784_out0 = v$G1_4092_out0;
assign v$COUT_1008_out0 = v$G1_4316_out0;
assign v$MULTI$OUT_13607_out0 = v$MULTI$REGIN_2870_out0;
assign v$MULTI$OUT_13608_out0 = v$MULTI$REGIN_2871_out0;
assign v$MULTI$OUT_1669_out0 = v$MULTI$OUT_13607_out0;
assign v$MULTI$OUT_1670_out0 = v$MULTI$OUT_13608_out0;
assign v$CIN_9911_out0 = v$COUT_784_out0;
assign v$CIN_10135_out0 = v$COUT_1008_out0;
assign v$RD_6077_out0 = v$CIN_9911_out0;
assign v$RD_6541_out0 = v$CIN_10135_out0;
assign v$G1_7932_out0 = ((v$RD_6077_out0 && !v$RM_11517_out0) || (!v$RD_6077_out0) && v$RM_11517_out0);
assign v$G1_8396_out0 = ((v$RD_6541_out0 && !v$RM_11981_out0) || (!v$RD_6541_out0) && v$RM_11981_out0);
assign v$G2_12468_out0 = v$RD_6077_out0 && v$RM_11517_out0;
assign v$G2_12932_out0 = v$RD_6541_out0 && v$RM_11981_out0;
assign v$CARRY_5077_out0 = v$G2_12468_out0;
assign v$CARRY_5541_out0 = v$G2_12932_out0;
assign v$S_9078_out0 = v$G1_7932_out0;
assign v$S_9542_out0 = v$G1_8396_out0;
assign v$S_1322_out0 = v$S_9078_out0;
assign v$S_1546_out0 = v$S_9542_out0;
assign v$G1_4098_out0 = v$CARRY_5077_out0 || v$CARRY_5076_out0;
assign v$G1_4322_out0 = v$CARRY_5541_out0 || v$CARRY_5540_out0;
assign v$COUT_790_out0 = v$G1_4098_out0;
assign v$COUT_1014_out0 = v$G1_4322_out0;
assign v$_4788_out0 = { v$S_1316_out0,v$S_1322_out0 };
assign v$_4803_out0 = { v$S_1540_out0,v$S_1546_out0 };
assign v$CIN_9906_out0 = v$COUT_790_out0;
assign v$CIN_10130_out0 = v$COUT_1014_out0;
assign v$RD_6067_out0 = v$CIN_9906_out0;
assign v$RD_6531_out0 = v$CIN_10130_out0;
assign v$G1_7922_out0 = ((v$RD_6067_out0 && !v$RM_11507_out0) || (!v$RD_6067_out0) && v$RM_11507_out0);
assign v$G1_8386_out0 = ((v$RD_6531_out0 && !v$RM_11971_out0) || (!v$RD_6531_out0) && v$RM_11971_out0);
assign v$G2_12458_out0 = v$RD_6067_out0 && v$RM_11507_out0;
assign v$G2_12922_out0 = v$RD_6531_out0 && v$RM_11971_out0;
assign v$CARRY_5067_out0 = v$G2_12458_out0;
assign v$CARRY_5531_out0 = v$G2_12922_out0;
assign v$S_9068_out0 = v$G1_7922_out0;
assign v$S_9532_out0 = v$G1_8386_out0;
assign v$S_1317_out0 = v$S_9068_out0;
assign v$S_1541_out0 = v$S_9532_out0;
assign v$G1_4093_out0 = v$CARRY_5067_out0 || v$CARRY_5066_out0;
assign v$G1_4317_out0 = v$CARRY_5531_out0 || v$CARRY_5530_out0;
assign v$COUT_785_out0 = v$G1_4093_out0;
assign v$COUT_1009_out0 = v$G1_4317_out0;
assign v$_2558_out0 = { v$_4788_out0,v$S_1317_out0 };
assign v$_2573_out0 = { v$_4803_out0,v$S_1541_out0 };
assign v$CIN_9901_out0 = v$COUT_785_out0;
assign v$CIN_10125_out0 = v$COUT_1009_out0;
assign v$RD_6056_out0 = v$CIN_9901_out0;
assign v$RD_6520_out0 = v$CIN_10125_out0;
assign v$G1_7911_out0 = ((v$RD_6056_out0 && !v$RM_11496_out0) || (!v$RD_6056_out0) && v$RM_11496_out0);
assign v$G1_8375_out0 = ((v$RD_6520_out0 && !v$RM_11960_out0) || (!v$RD_6520_out0) && v$RM_11960_out0);
assign v$G2_12447_out0 = v$RD_6056_out0 && v$RM_11496_out0;
assign v$G2_12911_out0 = v$RD_6520_out0 && v$RM_11960_out0;
assign v$CARRY_5056_out0 = v$G2_12447_out0;
assign v$CARRY_5520_out0 = v$G2_12911_out0;
assign v$S_9057_out0 = v$G1_7911_out0;
assign v$S_9521_out0 = v$G1_8375_out0;
assign v$S_1312_out0 = v$S_9057_out0;
assign v$S_1536_out0 = v$S_9521_out0;
assign v$G1_4088_out0 = v$CARRY_5056_out0 || v$CARRY_5055_out0;
assign v$G1_4312_out0 = v$CARRY_5520_out0 || v$CARRY_5519_out0;
assign v$COUT_780_out0 = v$G1_4088_out0;
assign v$COUT_1004_out0 = v$G1_4312_out0;
assign v$_7038_out0 = { v$_2558_out0,v$S_1312_out0 };
assign v$_7053_out0 = { v$_2573_out0,v$S_1536_out0 };
assign v$CIN_9900_out0 = v$COUT_780_out0;
assign v$CIN_10124_out0 = v$COUT_1004_out0;
assign v$RD_6054_out0 = v$CIN_9900_out0;
assign v$RD_6518_out0 = v$CIN_10124_out0;
assign v$G1_7909_out0 = ((v$RD_6054_out0 && !v$RM_11494_out0) || (!v$RD_6054_out0) && v$RM_11494_out0);
assign v$G1_8373_out0 = ((v$RD_6518_out0 && !v$RM_11958_out0) || (!v$RD_6518_out0) && v$RM_11958_out0);
assign v$G2_12445_out0 = v$RD_6054_out0 && v$RM_11494_out0;
assign v$G2_12909_out0 = v$RD_6518_out0 && v$RM_11958_out0;
assign v$CARRY_5054_out0 = v$G2_12445_out0;
assign v$CARRY_5518_out0 = v$G2_12909_out0;
assign v$S_9055_out0 = v$G1_7909_out0;
assign v$S_9519_out0 = v$G1_8373_out0;
assign v$S_1311_out0 = v$S_9055_out0;
assign v$S_1535_out0 = v$S_9519_out0;
assign v$G1_4087_out0 = v$CARRY_5054_out0 || v$CARRY_5053_out0;
assign v$G1_4311_out0 = v$CARRY_5518_out0 || v$CARRY_5517_out0;
assign v$COUT_779_out0 = v$G1_4087_out0;
assign v$COUT_1003_out0 = v$G1_4311_out0;
assign v$_13524_out0 = { v$_7038_out0,v$S_1311_out0 };
assign v$_13539_out0 = { v$_7053_out0,v$S_1535_out0 };
assign v$CIN_9907_out0 = v$COUT_779_out0;
assign v$CIN_10131_out0 = v$COUT_1003_out0;
assign v$RD_6069_out0 = v$CIN_9907_out0;
assign v$RD_6533_out0 = v$CIN_10131_out0;
assign v$G1_7924_out0 = ((v$RD_6069_out0 && !v$RM_11509_out0) || (!v$RD_6069_out0) && v$RM_11509_out0);
assign v$G1_8388_out0 = ((v$RD_6533_out0 && !v$RM_11973_out0) || (!v$RD_6533_out0) && v$RM_11973_out0);
assign v$G2_12460_out0 = v$RD_6069_out0 && v$RM_11509_out0;
assign v$G2_12924_out0 = v$RD_6533_out0 && v$RM_11973_out0;
assign v$CARRY_5069_out0 = v$G2_12460_out0;
assign v$CARRY_5533_out0 = v$G2_12924_out0;
assign v$S_9070_out0 = v$G1_7924_out0;
assign v$S_9534_out0 = v$G1_8388_out0;
assign v$S_1318_out0 = v$S_9070_out0;
assign v$S_1542_out0 = v$S_9534_out0;
assign v$G1_4094_out0 = v$CARRY_5069_out0 || v$CARRY_5068_out0;
assign v$G1_4318_out0 = v$CARRY_5533_out0 || v$CARRY_5532_out0;
assign v$COUT_786_out0 = v$G1_4094_out0;
assign v$COUT_1010_out0 = v$G1_4318_out0;
assign v$_3317_out0 = { v$_13524_out0,v$S_1318_out0 };
assign v$_3332_out0 = { v$_13539_out0,v$S_1542_out0 };
assign v$CIN_9908_out0 = v$COUT_786_out0;
assign v$CIN_10132_out0 = v$COUT_1010_out0;
assign v$RD_6071_out0 = v$CIN_9908_out0;
assign v$RD_6535_out0 = v$CIN_10132_out0;
assign v$G1_7926_out0 = ((v$RD_6071_out0 && !v$RM_11511_out0) || (!v$RD_6071_out0) && v$RM_11511_out0);
assign v$G1_8390_out0 = ((v$RD_6535_out0 && !v$RM_11975_out0) || (!v$RD_6535_out0) && v$RM_11975_out0);
assign v$G2_12462_out0 = v$RD_6071_out0 && v$RM_11511_out0;
assign v$G2_12926_out0 = v$RD_6535_out0 && v$RM_11975_out0;
assign v$CARRY_5071_out0 = v$G2_12462_out0;
assign v$CARRY_5535_out0 = v$G2_12926_out0;
assign v$S_9072_out0 = v$G1_7926_out0;
assign v$S_9536_out0 = v$G1_8390_out0;
assign v$S_1319_out0 = v$S_9072_out0;
assign v$S_1543_out0 = v$S_9536_out0;
assign v$G1_4095_out0 = v$CARRY_5071_out0 || v$CARRY_5070_out0;
assign v$G1_4319_out0 = v$CARRY_5535_out0 || v$CARRY_5534_out0;
assign v$COUT_787_out0 = v$G1_4095_out0;
assign v$COUT_1011_out0 = v$G1_4319_out0;
assign v$_7153_out0 = { v$_3317_out0,v$S_1319_out0 };
assign v$_7168_out0 = { v$_3332_out0,v$S_1543_out0 };
assign v$CIN_9910_out0 = v$COUT_787_out0;
assign v$CIN_10134_out0 = v$COUT_1011_out0;
assign v$RD_6075_out0 = v$CIN_9910_out0;
assign v$RD_6539_out0 = v$CIN_10134_out0;
assign v$G1_7930_out0 = ((v$RD_6075_out0 && !v$RM_11515_out0) || (!v$RD_6075_out0) && v$RM_11515_out0);
assign v$G1_8394_out0 = ((v$RD_6539_out0 && !v$RM_11979_out0) || (!v$RD_6539_out0) && v$RM_11979_out0);
assign v$G2_12466_out0 = v$RD_6075_out0 && v$RM_11515_out0;
assign v$G2_12930_out0 = v$RD_6539_out0 && v$RM_11979_out0;
assign v$CARRY_5075_out0 = v$G2_12466_out0;
assign v$CARRY_5539_out0 = v$G2_12930_out0;
assign v$S_9076_out0 = v$G1_7930_out0;
assign v$S_9540_out0 = v$G1_8394_out0;
assign v$S_1321_out0 = v$S_9076_out0;
assign v$S_1545_out0 = v$S_9540_out0;
assign v$G1_4097_out0 = v$CARRY_5075_out0 || v$CARRY_5074_out0;
assign v$G1_4321_out0 = v$CARRY_5539_out0 || v$CARRY_5538_out0;
assign v$COUT_789_out0 = v$G1_4097_out0;
assign v$COUT_1013_out0 = v$G1_4321_out0;
assign v$_4755_out0 = { v$_7153_out0,v$S_1321_out0 };
assign v$_4770_out0 = { v$_7168_out0,v$S_1545_out0 };
assign v$CIN_9903_out0 = v$COUT_789_out0;
assign v$CIN_10127_out0 = v$COUT_1013_out0;
assign v$RD_6061_out0 = v$CIN_9903_out0;
assign v$RD_6525_out0 = v$CIN_10127_out0;
assign v$G1_7916_out0 = ((v$RD_6061_out0 && !v$RM_11501_out0) || (!v$RD_6061_out0) && v$RM_11501_out0);
assign v$G1_8380_out0 = ((v$RD_6525_out0 && !v$RM_11965_out0) || (!v$RD_6525_out0) && v$RM_11965_out0);
assign v$G2_12452_out0 = v$RD_6061_out0 && v$RM_11501_out0;
assign v$G2_12916_out0 = v$RD_6525_out0 && v$RM_11965_out0;
assign v$CARRY_5061_out0 = v$G2_12452_out0;
assign v$CARRY_5525_out0 = v$G2_12916_out0;
assign v$S_9062_out0 = v$G1_7916_out0;
assign v$S_9526_out0 = v$G1_8380_out0;
assign v$S_1314_out0 = v$S_9062_out0;
assign v$S_1538_out0 = v$S_9526_out0;
assign v$G1_4090_out0 = v$CARRY_5061_out0 || v$CARRY_5060_out0;
assign v$G1_4314_out0 = v$CARRY_5525_out0 || v$CARRY_5524_out0;
assign v$COUT_782_out0 = v$G1_4090_out0;
assign v$COUT_1006_out0 = v$G1_4314_out0;
assign v$_6932_out0 = { v$_4755_out0,v$S_1314_out0 };
assign v$_6947_out0 = { v$_4770_out0,v$S_1538_out0 };
assign v$CIN_9904_out0 = v$COUT_782_out0;
assign v$CIN_10128_out0 = v$COUT_1006_out0;
assign v$RD_6063_out0 = v$CIN_9904_out0;
assign v$RD_6527_out0 = v$CIN_10128_out0;
assign v$G1_7918_out0 = ((v$RD_6063_out0 && !v$RM_11503_out0) || (!v$RD_6063_out0) && v$RM_11503_out0);
assign v$G1_8382_out0 = ((v$RD_6527_out0 && !v$RM_11967_out0) || (!v$RD_6527_out0) && v$RM_11967_out0);
assign v$G2_12454_out0 = v$RD_6063_out0 && v$RM_11503_out0;
assign v$G2_12918_out0 = v$RD_6527_out0 && v$RM_11967_out0;
assign v$CARRY_5063_out0 = v$G2_12454_out0;
assign v$CARRY_5527_out0 = v$G2_12918_out0;
assign v$S_9064_out0 = v$G1_7918_out0;
assign v$S_9528_out0 = v$G1_8382_out0;
assign v$S_1315_out0 = v$S_9064_out0;
assign v$S_1539_out0 = v$S_9528_out0;
assign v$G1_4091_out0 = v$CARRY_5063_out0 || v$CARRY_5062_out0;
assign v$G1_4315_out0 = v$CARRY_5527_out0 || v$CARRY_5526_out0;
assign v$COUT_783_out0 = v$G1_4091_out0;
assign v$COUT_1007_out0 = v$G1_4315_out0;
assign v$_5808_out0 = { v$_6932_out0,v$S_1315_out0 };
assign v$_5823_out0 = { v$_6947_out0,v$S_1539_out0 };
assign v$CIN_9909_out0 = v$COUT_783_out0;
assign v$CIN_10133_out0 = v$COUT_1007_out0;
assign v$RD_6073_out0 = v$CIN_9909_out0;
assign v$RD_6537_out0 = v$CIN_10133_out0;
assign v$G1_7928_out0 = ((v$RD_6073_out0 && !v$RM_11513_out0) || (!v$RD_6073_out0) && v$RM_11513_out0);
assign v$G1_8392_out0 = ((v$RD_6537_out0 && !v$RM_11977_out0) || (!v$RD_6537_out0) && v$RM_11977_out0);
assign v$G2_12464_out0 = v$RD_6073_out0 && v$RM_11513_out0;
assign v$G2_12928_out0 = v$RD_6537_out0 && v$RM_11977_out0;
assign v$CARRY_5073_out0 = v$G2_12464_out0;
assign v$CARRY_5537_out0 = v$G2_12928_out0;
assign v$S_9074_out0 = v$G1_7928_out0;
assign v$S_9538_out0 = v$G1_8392_out0;
assign v$S_1320_out0 = v$S_9074_out0;
assign v$S_1544_out0 = v$S_9538_out0;
assign v$G1_4096_out0 = v$CARRY_5073_out0 || v$CARRY_5072_out0;
assign v$G1_4320_out0 = v$CARRY_5537_out0 || v$CARRY_5536_out0;
assign v$COUT_788_out0 = v$G1_4096_out0;
assign v$COUT_1012_out0 = v$G1_4320_out0;
assign v$_2032_out0 = { v$_5808_out0,v$S_1320_out0 };
assign v$_2047_out0 = { v$_5823_out0,v$S_1544_out0 };
assign v$CIN_9897_out0 = v$COUT_788_out0;
assign v$CIN_10121_out0 = v$COUT_1012_out0;
assign v$RD_6048_out0 = v$CIN_9897_out0;
assign v$RD_6512_out0 = v$CIN_10121_out0;
assign v$G1_7903_out0 = ((v$RD_6048_out0 && !v$RM_11488_out0) || (!v$RD_6048_out0) && v$RM_11488_out0);
assign v$G1_8367_out0 = ((v$RD_6512_out0 && !v$RM_11952_out0) || (!v$RD_6512_out0) && v$RM_11952_out0);
assign v$G2_12439_out0 = v$RD_6048_out0 && v$RM_11488_out0;
assign v$G2_12903_out0 = v$RD_6512_out0 && v$RM_11952_out0;
assign v$CARRY_5048_out0 = v$G2_12439_out0;
assign v$CARRY_5512_out0 = v$G2_12903_out0;
assign v$S_9049_out0 = v$G1_7903_out0;
assign v$S_9513_out0 = v$G1_8367_out0;
assign v$S_1308_out0 = v$S_9049_out0;
assign v$S_1532_out0 = v$S_9513_out0;
assign v$G1_4084_out0 = v$CARRY_5048_out0 || v$CARRY_5047_out0;
assign v$G1_4308_out0 = v$CARRY_5512_out0 || v$CARRY_5511_out0;
assign v$COUT_776_out0 = v$G1_4084_out0;
assign v$COUT_1000_out0 = v$G1_4308_out0;
assign v$_2799_out0 = { v$_2032_out0,v$S_1308_out0 };
assign v$_2814_out0 = { v$_2047_out0,v$S_1532_out0 };
assign v$CIN_9902_out0 = v$COUT_776_out0;
assign v$CIN_10126_out0 = v$COUT_1000_out0;
assign v$RD_6058_out0 = v$CIN_9902_out0;
assign v$RD_6522_out0 = v$CIN_10126_out0;
assign v$G1_7913_out0 = ((v$RD_6058_out0 && !v$RM_11498_out0) || (!v$RD_6058_out0) && v$RM_11498_out0);
assign v$G1_8377_out0 = ((v$RD_6522_out0 && !v$RM_11962_out0) || (!v$RD_6522_out0) && v$RM_11962_out0);
assign v$G2_12449_out0 = v$RD_6058_out0 && v$RM_11498_out0;
assign v$G2_12913_out0 = v$RD_6522_out0 && v$RM_11962_out0;
assign v$CARRY_5058_out0 = v$G2_12449_out0;
assign v$CARRY_5522_out0 = v$G2_12913_out0;
assign v$S_9059_out0 = v$G1_7913_out0;
assign v$S_9523_out0 = v$G1_8377_out0;
assign v$S_1313_out0 = v$S_9059_out0;
assign v$S_1537_out0 = v$S_9523_out0;
assign v$G1_4089_out0 = v$CARRY_5058_out0 || v$CARRY_5057_out0;
assign v$G1_4313_out0 = v$CARRY_5522_out0 || v$CARRY_5521_out0;
assign v$COUT_781_out0 = v$G1_4089_out0;
assign v$COUT_1005_out0 = v$G1_4313_out0;
assign v$_1831_out0 = { v$_2799_out0,v$S_1313_out0 };
assign v$_1846_out0 = { v$_2814_out0,v$S_1537_out0 };
assign v$CIN_9898_out0 = v$COUT_781_out0;
assign v$CIN_10122_out0 = v$COUT_1005_out0;
assign v$RD_6050_out0 = v$CIN_9898_out0;
assign v$RD_6514_out0 = v$CIN_10122_out0;
assign v$G1_7905_out0 = ((v$RD_6050_out0 && !v$RM_11490_out0) || (!v$RD_6050_out0) && v$RM_11490_out0);
assign v$G1_8369_out0 = ((v$RD_6514_out0 && !v$RM_11954_out0) || (!v$RD_6514_out0) && v$RM_11954_out0);
assign v$G2_12441_out0 = v$RD_6050_out0 && v$RM_11490_out0;
assign v$G2_12905_out0 = v$RD_6514_out0 && v$RM_11954_out0;
assign v$CARRY_5050_out0 = v$G2_12441_out0;
assign v$CARRY_5514_out0 = v$G2_12905_out0;
assign v$S_9051_out0 = v$G1_7905_out0;
assign v$S_9515_out0 = v$G1_8369_out0;
assign v$S_1309_out0 = v$S_9051_out0;
assign v$S_1533_out0 = v$S_9515_out0;
assign v$G1_4085_out0 = v$CARRY_5050_out0 || v$CARRY_5049_out0;
assign v$G1_4309_out0 = v$CARRY_5514_out0 || v$CARRY_5513_out0;
assign v$COUT_777_out0 = v$G1_4085_out0;
assign v$COUT_1001_out0 = v$G1_4309_out0;
assign v$_4555_out0 = { v$_1831_out0,v$S_1309_out0 };
assign v$_4570_out0 = { v$_1846_out0,v$S_1533_out0 };
assign v$RM_3446_out0 = v$COUT_777_out0;
assign v$RM_3670_out0 = v$COUT_1001_out0;
assign v$RM_11491_out0 = v$RM_3446_out0;
assign v$RM_11955_out0 = v$RM_3670_out0;
assign v$G1_7906_out0 = ((v$RD_6051_out0 && !v$RM_11491_out0) || (!v$RD_6051_out0) && v$RM_11491_out0);
assign v$G1_8370_out0 = ((v$RD_6515_out0 && !v$RM_11955_out0) || (!v$RD_6515_out0) && v$RM_11955_out0);
assign v$G2_12442_out0 = v$RD_6051_out0 && v$RM_11491_out0;
assign v$G2_12906_out0 = v$RD_6515_out0 && v$RM_11955_out0;
assign v$CARRY_5051_out0 = v$G2_12442_out0;
assign v$CARRY_5515_out0 = v$G2_12906_out0;
assign v$S_9052_out0 = v$G1_7906_out0;
assign v$S_9516_out0 = v$G1_8370_out0;
assign v$RM_11492_out0 = v$S_9052_out0;
assign v$RM_11956_out0 = v$S_9516_out0;
assign v$G1_7907_out0 = ((v$RD_6052_out0 && !v$RM_11492_out0) || (!v$RD_6052_out0) && v$RM_11492_out0);
assign v$G1_8371_out0 = ((v$RD_6516_out0 && !v$RM_11956_out0) || (!v$RD_6516_out0) && v$RM_11956_out0);
assign v$G2_12443_out0 = v$RD_6052_out0 && v$RM_11492_out0;
assign v$G2_12907_out0 = v$RD_6516_out0 && v$RM_11956_out0;
assign v$CARRY_5052_out0 = v$G2_12443_out0;
assign v$CARRY_5516_out0 = v$G2_12907_out0;
assign v$S_9053_out0 = v$G1_7907_out0;
assign v$S_9517_out0 = v$G1_8371_out0;
assign v$S_1310_out0 = v$S_9053_out0;
assign v$S_1534_out0 = v$S_9517_out0;
assign v$G1_4086_out0 = v$CARRY_5052_out0 || v$CARRY_5051_out0;
assign v$G1_4310_out0 = v$CARRY_5516_out0 || v$CARRY_5515_out0;
assign v$COUT_778_out0 = v$G1_4086_out0;
assign v$COUT_1002_out0 = v$G1_4310_out0;
assign v$_10657_out0 = { v$_4555_out0,v$S_1310_out0 };
assign v$_10672_out0 = { v$_4570_out0,v$S_1534_out0 };
assign v$_10952_out0 = { v$_10657_out0,v$COUT_778_out0 };
assign v$_10967_out0 = { v$_10672_out0,v$COUT_1002_out0 };
assign v$COUT_10922_out0 = v$_10952_out0;
assign v$COUT_10937_out0 = v$_10967_out0;
assign v$_212_out0 = { v$_403_out0,v$COUT_10922_out0 };
assign v$_213_out0 = { v$_404_out0,v$COUT_10937_out0 };
assign v$FLOATING$MULTI_7697_out0 = v$_212_out0;
assign v$FLOATING$MULTI_7698_out0 = v$_213_out0;
assign v$32BIT$MULTI_1183_out0 = v$FLOATING$MULTI_7697_out0;
assign v$32BIT$MULTI_1184_out0 = v$FLOATING$MULTI_7698_out0;
assign v$32BITPRODUCT_82_out0 = v$32BIT$MULTI_1183_out0;
assign v$32BITPRODUCT_83_out0 = v$32BIT$MULTI_1184_out0;
assign v$32BITPRODUCT_12249_out0 = v$32BITPRODUCT_82_out0;
assign v$32BITPRODUCT_12250_out0 = v$32BITPRODUCT_83_out0;
assign v$SEL7_4850_out0 = v$32BITPRODUCT_12249_out0[21:10];
assign v$SEL7_4851_out0 = v$32BITPRODUCT_12250_out0[21:10];
assign v$MULTI$PRODUCT_7104_out0 = v$SEL7_4850_out0;
assign v$MULTI$PRODUCT_7105_out0 = v$SEL7_4851_out0;
assign v$MUX8_13785_out0 = v$MULTI$INSTRUCTION_2451_out0 ? v$MULTI$PRODUCT_7104_out0 : v$SEL8_10686_out0;
assign v$MUX8_13786_out0 = v$MULTI$INSTRUCTION_2452_out0 ? v$MULTI$PRODUCT_7105_out0 : v$SEL8_10687_out0;
assign v$SEL3_1143_out0 = v$MUX8_13785_out0[11:11];
assign v$SEL3_1144_out0 = v$MUX8_13786_out0[11:11];
assign v$SEL5_3049_out0 = v$MUX8_13785_out0[10:10];
assign v$SEL5_3050_out0 = v$MUX8_13786_out0[10:10];
assign v$SEL2_13496_out0 = v$MUX8_13785_out0[10:0];
assign v$SEL2_13497_out0 = v$MUX8_13786_out0[10:0];
assign v$SEL6_3991_out0 = v$SEL2_13496_out0[8:0];
assign v$SEL6_3992_out0 = v$SEL2_13497_out0[8:0];
assign v$BIT10_7009_out0 = v$SEL5_3049_out0;
assign v$BIT10_7010_out0 = v$SEL5_3050_out0;
assign v$OVERFLOW_10492_out0 = v$SEL3_1143_out0;
assign v$OVERFLOW_10493_out0 = v$SEL3_1144_out0;
assign v$SEL4_11225_out0 = v$SEL2_13496_out0[9:0];
assign v$SEL4_11226_out0 = v$SEL2_13497_out0[9:0];
assign v$SEL9_13753_out0 = v$SEL2_13496_out0[10:1];
assign v$SEL9_13754_out0 = v$SEL2_13497_out0[10:1];
assign v$G3_2690_out0 = v$BIT10_7009_out0 || v$OVERFLOW_10492_out0;
assign v$G3_2691_out0 = v$BIT10_7010_out0 || v$OVERFLOW_10493_out0;
assign v$_8677_out0 = { v$C9_3029_out0,v$SEL6_3991_out0 };
assign v$_8678_out0 = { v$C9_3030_out0,v$SEL6_3992_out0 };
assign v$MUX5_10260_out0 = v$SUBNORMAL_8808_out0 ? v$BIT10_7009_out0 : v$OVERFLOW_10492_out0;
assign v$MUX5_10261_out0 = v$SUBNORMAL_8809_out0 ? v$BIT10_7010_out0 : v$OVERFLOW_10493_out0;
assign v$MUX4_10357_out0 = v$OVERFLOW_10492_out0 ? v$SEL9_13753_out0 : v$SEL4_11225_out0;
assign v$MUX4_10358_out0 = v$OVERFLOW_10493_out0 ? v$SEL9_13754_out0 : v$SEL4_11226_out0;
assign v$G2_5840_out0 = !(v$G3_2690_out0 || v$SUBNORMAL_8808_out0);
assign v$G2_5841_out0 = !(v$G3_2691_out0 || v$SUBNORMAL_8809_out0);
assign v$UNDERFLOW_6916_out0 = v$G2_5840_out0;
assign v$UNDERFLOW_6917_out0 = v$G2_5841_out0;
assign v$G4_3235_out0 = v$UNDERFLOW_6916_out0 && v$G5_638_out0;
assign v$G4_3236_out0 = v$UNDERFLOW_6917_out0 && v$G5_639_out0;
assign v$MUX7_4481_out0 = v$UNDERFLOW_6916_out0 ? v$C10_11248_out0 : v$C8_2758_out0;
assign v$MUX7_4482_out0 = v$UNDERFLOW_6917_out0 ? v$C10_11249_out0 : v$C8_2759_out0;
assign {v$A7_2719_out1,v$A7_2719_out0 } = v$EXP_2441_out0 + v$MUX7_4481_out0 + v$MUX5_10260_out0;
assign {v$A7_2720_out1,v$A7_2720_out0 } = v$EXP_2442_out0 + v$MUX7_4482_out0 + v$MUX5_10261_out0;
assign v$MUX6_10350_out0 = v$G4_3235_out0 ? v$_8677_out0 : v$MUX4_10357_out0;
assign v$MUX6_10351_out0 = v$G4_3236_out0 ? v$_8678_out0 : v$MUX4_10358_out0;
assign v$SIG$ANS_439_out0 = v$MUX6_10350_out0;
assign v$SIG$ANS_440_out0 = v$MUX6_10351_out0;
assign v$NOTUSED3_10550_out0 = v$A7_2719_out1;
assign v$NOTUSED3_10551_out0 = v$A7_2720_out1;
assign v$EXP$ANS_13748_out0 = v$A7_2719_out0;
assign v$EXP$ANS_13749_out0 = v$A7_2720_out0;
assign v$EXP$ANS_2008_out0 = v$EXP$ANS_13748_out0;
assign v$EXP$ANS_2009_out0 = v$EXP$ANS_13749_out0;
assign v$SIG$ANS_2335_out0 = v$SIG$ANS_439_out0;
assign v$SIG$ANS_2336_out0 = v$SIG$ANS_440_out0;
assign v$_2610_out0 = { v$EXP$ANS_2008_out0,v$SIGN$ANS_8650_out0 };
assign v$_2611_out0 = { v$EXP$ANS_2009_out0,v$SIGN$ANS_8651_out0 };
assign v$SIG$ANS_3276_out0 = v$SIG$ANS_2335_out0;
assign v$SIG$ANS_3277_out0 = v$SIG$ANS_2336_out0;
assign v$EXP$ANS_10487_out0 = v$EXP$ANS_2008_out0;
assign v$EXP$ANS_10488_out0 = v$EXP$ANS_2009_out0;
assign v$SIG$ANS_10296_out0 = v$SIG$ANS_3276_out0;
assign v$SIG$ANS_10297_out0 = v$SIG$ANS_3277_out0;
assign v$_10449_out0 = { v$SIG$ANS_2335_out0,v$_2610_out0 };
assign v$_10450_out0 = { v$SIG$ANS_2336_out0,v$_2611_out0 };
assign v$EXP$ANS_11059_out0 = v$EXP$ANS_10487_out0;
assign v$EXP$ANS_11060_out0 = v$EXP$ANS_10488_out0;
assign v$16BIT$WORD$ANSWER_8821_out0 = v$_10449_out0;
assign v$16BIT$WORD$ANSWER_8822_out0 = v$_10450_out0;
assign v$FLOATING$REGISTER$IN_562_out0 = v$16BIT$WORD$ANSWER_8821_out0;
assign v$FLOATING$REGISTER$IN_563_out0 = v$16BIT$WORD$ANSWER_8822_out0;
assign v$MUX12_1714_out0 = v$FLOATING$EN$ALU_634_out0 ? v$FLOATING$REGISTER$IN_562_out0 : v$ALUOUT_4607_out0;
assign v$MUX12_1715_out0 = v$FLOATING$EN$ALU_635_out0 ? v$FLOATING$REGISTER$IN_563_out0 : v$ALUOUT_4608_out0;
assign v$MUX5_2606_out0 = v$FLOATING$INS_13797_out0 ? v$FLOATING$REGISTER$IN_562_out0 : v$MULTI$REGIN_2870_out0;
assign v$MUX5_2607_out0 = v$FLOATING$INS_13798_out0 ? v$FLOATING$REGISTER$IN_563_out0 : v$MULTI$REGIN_2871_out0;
assign v$MUX4_10_out0 = v$MULTI$OPCODE_3020_out0 ? v$MUX5_2606_out0 : v$LS$REGIN_3303_out0;
assign v$MUX4_11_out0 = v$MULTI$OPCODE_3021_out0 ? v$MUX5_2607_out0 : v$LS$REGIN_3304_out0;
assign v$MUX11_13745_out0 = v$IR15_2464_out0 ? v$MUX12_1714_out0 : v$MUX4_10_out0;
assign v$MUX11_13746_out0 = v$IR15_2465_out0 ? v$MUX12_1715_out0 : v$MUX4_11_out0;
assign v$DIN_2266_out0 = v$MUX11_13745_out0;
assign v$DIN_2267_out0 = v$MUX11_13746_out0;
assign v$DIN3_10310_out0 = v$MUX11_13745_out0;
assign v$DIN3_10311_out0 = v$MUX11_13746_out0;
assign v$DIN_9798_out0 = v$DIN_2266_out0;
assign v$DIN_9799_out0 = v$DIN_2267_out0;


endmodule
